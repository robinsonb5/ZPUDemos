-- ZPU
--
-- Copyright 2004-2008 oharboe - �yvind Harboe - oyvind.harboe@zylin.com
-- Modified by Alastair M. Robinson for the ZPUFlex project.
--
-- The FreeBSD license
-- 
-- Redistribution and use in source and binary forms, with or without
-- modification, are permitted provided that the following conditions
-- are met:
-- 
-- 1. Redistributions of source code must retain the above copyright
--    notice, this list of conditions and the following disclaimer.
-- 2. Redistributions in binary form must reproduce the above
--    copyright notice, this list of conditions and the following
--    disclaimer in the documentation and/or other materials
--    provided with the distribution.
-- 
-- THIS SOFTWARE IS PROVIDED BY THE ZPU PROJECT ``AS IS'' AND ANY
-- EXPRESS OR IMPLIED WARRANTIES, INCLUDING, BUT NOT LIMITED TO,
-- THE IMPLIED WARRANTIES OF MERCHANTABILITY AND FITNESS FOR A
-- PARTICULAR PURPOSE ARE DISCLAIMED. IN NO EVENT SHALL THE
-- ZPU PROJECT OR CONTRIBUTORS BE LIABLE FOR ANY DIRECT,
-- INDIRECT, INCIDENTAL, SPECIAL, EXEMPLARY, OR CONSEQUENTIAL DAMAGES
-- (INCLUDING, BUT NOT LIMITED TO, PROCUREMENT OF SUBSTITUTE GOODS
-- OR SERVICES; LOSS OF USE, DATA, OR PROFITS; OR BUSINESS INTERRUPTION)
-- HOWEVER CAUSED AND ON ANY THEORY OF LIABILITY, WHETHER IN CONTRACT,
-- STRICT LIABILITY, OR TORT (INCLUDING NEGLIGENCE OR OTHERWISE)
-- ARISING IN ANY WAY OUT OF THE USE OF THIS SOFTWARE, EVEN IF
-- ADVISED OF THE POSSIBILITY OF SUCH DAMAGE.
-- 
-- The views and conclusions contained in the software and documentation
-- are those of the authors and should not be interpreted as representing
-- official policies, either expressed or implied, of the ZPU Project.

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;


library work;
use work.zpupkg.all;

entity SDBootstrap_ROM is
generic
	(
		maxAddrBitBRAM : integer := maxAddrBitBRAMLimit -- Specify your actual ROM size to save LEs and unnecessary block RAM usage.
	);
port (
	clk : in std_logic;
	areset : in std_logic := '0';
	from_zpu : in ZPU_ToROM;
	to_zpu : out ZPU_FromROM
);
end SDBootstrap_ROM;

architecture arch of SDBootstrap_ROM is

type ram_type is array(natural range 0 to ((2**(maxAddrBitBRAM+1))/4)-1) of std_logic_vector(wordSize-1 downto 0);

shared variable ram : ram_type :=
(
     0 => x"84808080",
     1 => x"8c0b8480",
     2 => x"8081e004",
     3 => x"00848080",
     4 => x"808c04ff",
     5 => x"0d800404",
     6 => x"40000017",
     7 => x"00000000",
     8 => x"0b83ffe0",
     9 => x"80080b83",
    10 => x"ffe08408",
    11 => x"0b83ffe0",
    12 => x"88088480",
    13 => x"80809808",
    14 => x"2d0b83ff",
    15 => x"e0880c0b",
    16 => x"83ffe084",
    17 => x"0c0b83ff",
    18 => x"e0800c04",
    19 => x"00000000",
    20 => x"00000000",
    21 => x"00000000",
    22 => x"00000000",
    23 => x"00000000",
    24 => x"71fd0608",
    25 => x"72830609",
    26 => x"81058205",
    27 => x"832b2a83",
    28 => x"ffff0652",
    29 => x"0471fc06",
    30 => x"08728306",
    31 => x"09810583",
    32 => x"05101010",
    33 => x"2a81ff06",
    34 => x"520471fd",
    35 => x"060883ff",
    36 => x"ff738306",
    37 => x"09810582",
    38 => x"05832b2b",
    39 => x"09067383",
    40 => x"ffff0673",
    41 => x"83060981",
    42 => x"05820583",
    43 => x"2b0b2b07",
    44 => x"72fc060c",
    45 => x"51510471",
    46 => x"fc060884",
    47 => x"8080ad98",
    48 => x"73830610",
    49 => x"10050806",
    50 => x"7381ff06",
    51 => x"73830609",
    52 => x"81058305",
    53 => x"1010102b",
    54 => x"0772fc06",
    55 => x"0c515104",
    56 => x"83ffe080",
    57 => x"7083fff6",
    58 => x"a8278e38",
    59 => x"80717084",
    60 => x"05530c84",
    61 => x"808081e4",
    62 => x"04848080",
    63 => x"808c5184",
    64 => x"80809b80",
    65 => x"0402ec05",
    66 => x"0d765380",
    67 => x"5572752e",
    68 => x"be388754",
    69 => x"729c2a73",
    70 => x"842b5452",
    71 => x"71802e83",
    72 => x"38815589",
    73 => x"72258a38",
    74 => x"b7125284",
    75 => x"808082b4",
    76 => x"04b01252",
    77 => x"74802e89",
    78 => x"38715184",
    79 => x"808085a1",
    80 => x"2dff1454",
    81 => x"738025cc",
    82 => x"38848080",
    83 => x"82d704b0",
    84 => x"51848080",
    85 => x"85a12d80",
    86 => x"0b83ffe0",
    87 => x"800c0294",
    88 => x"050d0402",
    89 => x"c0050d02",
    90 => x"80c40557",
    91 => x"80707870",
    92 => x"84055a08",
    93 => x"72415f5d",
    94 => x"587c7084",
    95 => x"055e085a",
    96 => x"805b7998",
    97 => x"2a7a882b",
    98 => x"5b567589",
    99 => x"38775f84",
   100 => x"80808595",
   101 => x"047d802e",
   102 => x"81d33880",
   103 => x"5e7580e4",
   104 => x"2e8a3875",
   105 => x"80f82e09",
   106 => x"81068938",
   107 => x"76841871",
   108 => x"085e5854",
   109 => x"7580e42e",
   110 => x"a6387580",
   111 => x"e4268e38",
   112 => x"7580e32e",
   113 => x"80d93884",
   114 => x"808084ad",
   115 => x"047580f3",
   116 => x"2eb53875",
   117 => x"80f82e8f",
   118 => x"38848080",
   119 => x"84ad048a",
   120 => x"53848080",
   121 => x"83e90490",
   122 => x"5383ffe0",
   123 => x"e0527b51",
   124 => x"84808082",
   125 => x"852d83ff",
   126 => x"e0800883",
   127 => x"ffe0e05a",
   128 => x"55848080",
   129 => x"84c60476",
   130 => x"84187108",
   131 => x"70545b58",
   132 => x"54848080",
   133 => x"85c52d80",
   134 => x"55848080",
   135 => x"84c60476",
   136 => x"84187108",
   137 => x"58585484",
   138 => x"808084fd",
   139 => x"04a55184",
   140 => x"808085a1",
   141 => x"2d755184",
   142 => x"808085a1",
   143 => x"2d821858",
   144 => x"84808085",
   145 => x"880474ff",
   146 => x"16565480",
   147 => x"7425b938",
   148 => x"78708105",
   149 => x"5a848080",
   150 => x"80f52d70",
   151 => x"52568480",
   152 => x"8085a12d",
   153 => x"81185884",
   154 => x"808084c6",
   155 => x"0475a52e",
   156 => x"09810689",
   157 => x"38815e84",
   158 => x"80808588",
   159 => x"04755184",
   160 => x"808085a1",
   161 => x"2d811858",
   162 => x"811b5b83",
   163 => x"7b25fdf2",
   164 => x"3875fde5",
   165 => x"387e83ff",
   166 => x"e0800c02",
   167 => x"80c0050d",
   168 => x"0402f805",
   169 => x"0d7352c0",
   170 => x"0870882a",
   171 => x"70810651",
   172 => x"51517080",
   173 => x"2ef13871",
   174 => x"c00c7183",
   175 => x"ffe0800c",
   176 => x"0288050d",
   177 => x"0402e805",
   178 => x"0d807857",
   179 => x"55757084",
   180 => x"05570853",
   181 => x"80547298",
   182 => x"2a73882b",
   183 => x"54527180",
   184 => x"2ea238c0",
   185 => x"0870882a",
   186 => x"70810651",
   187 => x"51517080",
   188 => x"2ef13871",
   189 => x"c00c8115",
   190 => x"81155555",
   191 => x"837425d6",
   192 => x"3871ca38",
   193 => x"7483ffe0",
   194 => x"800c0298",
   195 => x"050d0402",
   196 => x"f4050dd4",
   197 => x"5281ff72",
   198 => x"0c710853",
   199 => x"81ff720c",
   200 => x"72882b83",
   201 => x"fe800672",
   202 => x"087081ff",
   203 => x"06515253",
   204 => x"81ff720c",
   205 => x"72710788",
   206 => x"2b720870",
   207 => x"81ff0651",
   208 => x"525381ff",
   209 => x"720c7271",
   210 => x"07882b72",
   211 => x"087081ff",
   212 => x"06720783",
   213 => x"ffe0800c",
   214 => x"5253028c",
   215 => x"050d0402",
   216 => x"ec050d76",
   217 => x"787181ff",
   218 => x"06705584",
   219 => x"8080ada8",
   220 => x"54555555",
   221 => x"84808082",
   222 => x"e32d72d4",
   223 => x"0c83fff1",
   224 => x"a0088538",
   225 => x"73892b54",
   226 => x"73528480",
   227 => x"80adb451",
   228 => x"84808082",
   229 => x"e32d7398",
   230 => x"2ad40c73",
   231 => x"902a7081",
   232 => x"ff06d40c",
   233 => x"5373882a",
   234 => x"7081ff06",
   235 => x"d40c5373",
   236 => x"81ff06d4",
   237 => x"0c74902a",
   238 => x"7081ff06",
   239 => x"70548480",
   240 => x"80adc053",
   241 => x"51538480",
   242 => x"8082e32d",
   243 => x"72d40cd4",
   244 => x"087081ff",
   245 => x"06515382",
   246 => x"b8bf5472",
   247 => x"81ff2e09",
   248 => x"81069438",
   249 => x"81ff0bd4",
   250 => x"0cd40870",
   251 => x"81ff06ff",
   252 => x"16565153",
   253 => x"73e53872",
   254 => x"52848080",
   255 => x"add05184",
   256 => x"808082e3",
   257 => x"2d7283ff",
   258 => x"e0800c02",
   259 => x"94050d04",
   260 => x"02fc050d",
   261 => x"81c75181",
   262 => x"ff0bd40c",
   263 => x"ff115170",
   264 => x"8025f438",
   265 => x"0284050d",
   266 => x"0402f005",
   267 => x"0d848080",
   268 => x"88902d81",
   269 => x"9c9f5380",
   270 => x"5287fc80",
   271 => x"f7518480",
   272 => x"8086df2d",
   273 => x"83ffe080",
   274 => x"085483ff",
   275 => x"e0800881",
   276 => x"2e098106",
   277 => x"b43881ff",
   278 => x"0bd40c82",
   279 => x"0a52849c",
   280 => x"80e95184",
   281 => x"808086df",
   282 => x"2d83ffe0",
   283 => x"80088e38",
   284 => x"81ff0bd4",
   285 => x"0c735384",
   286 => x"808089a2",
   287 => x"04848080",
   288 => x"88902d84",
   289 => x"8080899b",
   290 => x"0483ffe0",
   291 => x"80085284",
   292 => x"8080add4",
   293 => x"51848080",
   294 => x"82e32dff",
   295 => x"135372ff",
   296 => x"96387283",
   297 => x"ffe0800c",
   298 => x"0290050d",
   299 => x"0402f405",
   300 => x"0d81ff0b",
   301 => x"d40c8480",
   302 => x"80ade051",
   303 => x"84808085",
   304 => x"c52d9353",
   305 => x"805287fc",
   306 => x"80c15184",
   307 => x"808086df",
   308 => x"2d83ffe0",
   309 => x"80088e38",
   310 => x"81ff0bd4",
   311 => x"0c815384",
   312 => x"80808a83",
   313 => x"0483ffe0",
   314 => x"80085284",
   315 => x"8080ade4",
   316 => x"51848080",
   317 => x"82e32d84",
   318 => x"80808890",
   319 => x"2dff1353",
   320 => x"72c23872",
   321 => x"83ffe080",
   322 => x"0c028c05",
   323 => x"0d0402f4",
   324 => x"050d8480",
   325 => x"8088902d",
   326 => x"83aa5284",
   327 => x"9c80c851",
   328 => x"84808086",
   329 => x"df2d83ff",
   330 => x"e0800883",
   331 => x"ffe08008",
   332 => x"53848080",
   333 => x"adf05253",
   334 => x"84808082",
   335 => x"e32d7281",
   336 => x"2ea13872",
   337 => x"52848080",
   338 => x"ae885184",
   339 => x"808082e3",
   340 => x"2d848080",
   341 => x"89ad2d84",
   342 => x"8080aea0",
   343 => x"51848080",
   344 => x"8b980484",
   345 => x"8080868f",
   346 => x"2d83ffe0",
   347 => x"800883ff",
   348 => x"ff065372",
   349 => x"83aa2e80",
   350 => x"d33883ff",
   351 => x"e0800852",
   352 => x"848080ae",
   353 => x"88518480",
   354 => x"8082e32d",
   355 => x"84808089",
   356 => x"ad2d8480",
   357 => x"80aea851",
   358 => x"84808085",
   359 => x"c52d8480",
   360 => x"808bc404",
   361 => x"848080ae",
   362 => x"b8518480",
   363 => x"8085c52d",
   364 => x"81538480",
   365 => x"808d8204",
   366 => x"848080ae",
   367 => x"c0518480",
   368 => x"8082e32d",
   369 => x"80538480",
   370 => x"808d8204",
   371 => x"81ff0bd4",
   372 => x"0c848080",
   373 => x"aedc5184",
   374 => x"808085c5",
   375 => x"2db15384",
   376 => x"808088a9",
   377 => x"2d83ffe0",
   378 => x"8008802e",
   379 => x"81873880",
   380 => x"5287fc80",
   381 => x"fa518480",
   382 => x"8086df2d",
   383 => x"83ffe080",
   384 => x"0880e038",
   385 => x"83ffe080",
   386 => x"08528480",
   387 => x"80aef451",
   388 => x"84808082",
   389 => x"e32d81ff",
   390 => x"0bd40cd4",
   391 => x"087081ff",
   392 => x"06705484",
   393 => x"8080af80",
   394 => x"53515384",
   395 => x"808082e3",
   396 => x"2d81ff0b",
   397 => x"d40c81ff",
   398 => x"0bd40c81",
   399 => x"ff0bd40c",
   400 => x"81ff0bd4",
   401 => x"0c72862a",
   402 => x"70810651",
   403 => x"5372fed4",
   404 => x"38848080",
   405 => x"af905184",
   406 => x"808085c5",
   407 => x"2d848080",
   408 => x"8d820483",
   409 => x"ffe08008",
   410 => x"52848080",
   411 => x"aef45184",
   412 => x"808082e3",
   413 => x"2d72822e",
   414 => x"febe38ff",
   415 => x"135372fe",
   416 => x"de387283",
   417 => x"ffe0800c",
   418 => x"028c050d",
   419 => x"0402e805",
   420 => x"0d785681",
   421 => x"ff0bd40c",
   422 => x"d008708f",
   423 => x"2a708106",
   424 => x"51515372",
   425 => x"f3388281",
   426 => x"0bd00c81",
   427 => x"ff0bd40c",
   428 => x"775287fc",
   429 => x"80d85184",
   430 => x"808086df",
   431 => x"2d83ffe0",
   432 => x"8008802e",
   433 => x"95388480",
   434 => x"80af9451",
   435 => x"84808085",
   436 => x"c52d8153",
   437 => x"8480808e",
   438 => x"d20481ff",
   439 => x"0bd40c81",
   440 => x"fe0bd40c",
   441 => x"80ff5575",
   442 => x"70840557",
   443 => x"0870982a",
   444 => x"d40c7090",
   445 => x"2c7081ff",
   446 => x"06d40c54",
   447 => x"70882c70",
   448 => x"81ff06d4",
   449 => x"0c547081",
   450 => x"ff06d40c",
   451 => x"54ff1555",
   452 => x"748025d3",
   453 => x"3881ff0b",
   454 => x"d40c81ff",
   455 => x"0bd40c81",
   456 => x"ff0bd40c",
   457 => x"868da054",
   458 => x"81ff0bd4",
   459 => x"0cd40881",
   460 => x"ff065574",
   461 => x"8738ff14",
   462 => x"5473ed38",
   463 => x"81ff0bd4",
   464 => x"0cd00870",
   465 => x"8f2a7081",
   466 => x"06515153",
   467 => x"72f33872",
   468 => x"d00c7283",
   469 => x"ffe0800c",
   470 => x"0298050d",
   471 => x"0402ec05",
   472 => x"0d767853",
   473 => x"54805580",
   474 => x"dbc6df53",
   475 => x"81ff0bd4",
   476 => x"0cd40870",
   477 => x"81ff0651",
   478 => x"517081fe",
   479 => x"2e098106",
   480 => x"80eb3880",
   481 => x"0b83fff1",
   482 => x"c40c8372",
   483 => x"25ab3884",
   484 => x"8080868f",
   485 => x"2d83ffe0",
   486 => x"80087470",
   487 => x"8405560c",
   488 => x"83fff1c4",
   489 => x"0883ffe0",
   490 => x"80080583",
   491 => x"fff1c40c",
   492 => x"fc125284",
   493 => x"80808f8a",
   494 => x"04807225",
   495 => x"a83881ff",
   496 => x"0bd40cff",
   497 => x"74708105",
   498 => x"56848080",
   499 => x"81b72d83",
   500 => x"fff1c408",
   501 => x"81ff0583",
   502 => x"fff1c40c",
   503 => x"ff125284",
   504 => x"80808fb9",
   505 => x"04815584",
   506 => x"80808ff4",
   507 => x"04ff1353",
   508 => x"72fef938",
   509 => x"81ff0bd4",
   510 => x"0c7483ff",
   511 => x"e0800c02",
   512 => x"94050d04",
   513 => x"02e0050d",
   514 => x"805287fc",
   515 => x"80c95184",
   516 => x"808086df",
   517 => x"2d83ffe0",
   518 => x"80085284",
   519 => x"8080afa4",
   520 => x"51848080",
   521 => x"82e32d92",
   522 => x"5283fff1",
   523 => x"b0518480",
   524 => x"808edd2d",
   525 => x"805583ff",
   526 => x"f1b01584",
   527 => x"808080f5",
   528 => x"2d528480",
   529 => x"80adb851",
   530 => x"84808082",
   531 => x"e32d8115",
   532 => x"55917525",
   533 => x"e1388480",
   534 => x"80addc51",
   535 => x"84808085",
   536 => x"c52d83ff",
   537 => x"f1b00b84",
   538 => x"808080f5",
   539 => x"2d81c006",
   540 => x"557480c0",
   541 => x"2e098106",
   542 => x"80c23883",
   543 => x"fff1b70b",
   544 => x"84808080",
   545 => x"f52d83ff",
   546 => x"f1b80b84",
   547 => x"808080f5",
   548 => x"2d71902b",
   549 => x"71882b07",
   550 => x"83fff1b9",
   551 => x"0b848080",
   552 => x"80f52d71",
   553 => x"81fffe80",
   554 => x"06077088",
   555 => x"80298880",
   556 => x"05515157",
   557 => x"59578480",
   558 => x"80938504",
   559 => x"83fff1b9",
   560 => x"0b848080",
   561 => x"80f52d70",
   562 => x"10860683",
   563 => x"fff1ba0b",
   564 => x"84808080",
   565 => x"f52d7087",
   566 => x"2a720783",
   567 => x"fff1b50b",
   568 => x"84808080",
   569 => x"f52d8f06",
   570 => x"83fff1b6",
   571 => x"0b848080",
   572 => x"80f52d70",
   573 => x"8a2b9880",
   574 => x"0683fff1",
   575 => x"b70b8480",
   576 => x"8080f52d",
   577 => x"70822b72",
   578 => x"0783fff1",
   579 => x"b80b8480",
   580 => x"8080f52d",
   581 => x"70862a72",
   582 => x"07705f76",
   583 => x"5e775d84",
   584 => x"8080afb8",
   585 => x"5c525252",
   586 => x"525c5354",
   587 => x"525a5657",
   588 => x"84808082",
   589 => x"e32d8215",
   590 => x"81712b70",
   591 => x"54848080",
   592 => x"afe85351",
   593 => x"55848080",
   594 => x"82e32d81",
   595 => x"772b7676",
   596 => x"29167155",
   597 => x"70548480",
   598 => x"80aff453",
   599 => x"56578480",
   600 => x"8082e32d",
   601 => x"84807725",
   602 => x"8e387410",
   603 => x"77812c58",
   604 => x"55848080",
   605 => x"92e40474",
   606 => x"52848080",
   607 => x"b08c5184",
   608 => x"808082e3",
   609 => x"2d7483ff",
   610 => x"e0800c02",
   611 => x"a0050d04",
   612 => x"02f0050d",
   613 => x"810b83ff",
   614 => x"f1a00c84",
   615 => x"8080b0a4",
   616 => x"51848080",
   617 => x"85c52d87",
   618 => x"54d00870",
   619 => x"8f2a7081",
   620 => x"06515153",
   621 => x"72f33872",
   622 => x"d00c8480",
   623 => x"8088902d",
   624 => x"848080b0",
   625 => x"a8518480",
   626 => x"8085c52d",
   627 => x"d008708f",
   628 => x"2a708106",
   629 => x"51515372",
   630 => x"f338810b",
   631 => x"d00c7252",
   632 => x"84d480c0",
   633 => x"51848080",
   634 => x"86df2d83",
   635 => x"ffe08008",
   636 => x"812e0981",
   637 => x"06873883",
   638 => x"ffe08008",
   639 => x"54848080",
   640 => x"b0b85184",
   641 => x"808085c5",
   642 => x"2d73822e",
   643 => x"bf38ff14",
   644 => x"5473ff95",
   645 => x"38848080",
   646 => x"b0cc5184",
   647 => x"808085c5",
   648 => x"2d848080",
   649 => x"8a8e2d83",
   650 => x"ffe08008",
   651 => x"83fff1a0",
   652 => x"0c83ffe0",
   653 => x"8008802e",
   654 => x"b1388480",
   655 => x"80b0e851",
   656 => x"84808085",
   657 => x"c52d8480",
   658 => x"80958304",
   659 => x"848080b0",
   660 => x"fc518480",
   661 => x"8085c52d",
   662 => x"848080b1",
   663 => x"84518480",
   664 => x"8085c52d",
   665 => x"84808095",
   666 => x"ce048480",
   667 => x"80b1a451",
   668 => x"84808085",
   669 => x"c52d8152",
   670 => x"87fc80d0",
   671 => x"51848080",
   672 => x"86df2d81",
   673 => x"ff0bd40c",
   674 => x"84808090",
   675 => x"842d83ff",
   676 => x"e0800883",
   677 => x"fff1a40c",
   678 => x"83ffe080",
   679 => x"08528480",
   680 => x"80b1c051",
   681 => x"84808082",
   682 => x"e32dd008",
   683 => x"708f2a70",
   684 => x"81065151",
   685 => x"5372f338",
   686 => x"72d00c81",
   687 => x"ff0bd40c",
   688 => x"848080b1",
   689 => x"d4518480",
   690 => x"8085c52d",
   691 => x"81537283",
   692 => x"ffe0800c",
   693 => x"0290050d",
   694 => x"0402e805",
   695 => x"0d775580",
   696 => x"5681ff0b",
   697 => x"d40cd008",
   698 => x"708f2a70",
   699 => x"81065151",
   700 => x"5473f338",
   701 => x"82810bd0",
   702 => x"0c81ff0b",
   703 => x"d40c7452",
   704 => x"87fc80d1",
   705 => x"51848080",
   706 => x"86df2d83",
   707 => x"ffe08008",
   708 => x"802e9b38",
   709 => x"83ffe080",
   710 => x"08537452",
   711 => x"848080b1",
   712 => x"e0518480",
   713 => x"8082e32d",
   714 => x"84808096",
   715 => x"d0048480",
   716 => x"52785184",
   717 => x"80808edd",
   718 => x"2d83ffe0",
   719 => x"800856d0",
   720 => x"08708f2a",
   721 => x"70810651",
   722 => x"515473f3",
   723 => x"3873d00c",
   724 => x"7583ffe0",
   725 => x"800c0298",
   726 => x"050d0402",
   727 => x"f4050d74",
   728 => x"70882a83",
   729 => x"fe800670",
   730 => x"72982a07",
   731 => x"72882b87",
   732 => x"fc808006",
   733 => x"71077398",
   734 => x"2b0783ff",
   735 => x"e0800c51",
   736 => x"5351028c",
   737 => x"050d0402",
   738 => x"f8050d02",
   739 => x"8e058480",
   740 => x"8080f52d",
   741 => x"74882b07",
   742 => x"7083ffff",
   743 => x"0683ffe0",
   744 => x"800c5102",
   745 => x"88050d04",
   746 => x"02f8050d",
   747 => x"7370902b",
   748 => x"71902a07",
   749 => x"83ffe080",
   750 => x"0c520288",
   751 => x"050d0402",
   752 => x"fc050d73",
   753 => x"81df06c9",
   754 => x"05517080",
   755 => x"258438a7",
   756 => x"11517284",
   757 => x"2b710783",
   758 => x"ffe0800c",
   759 => x"0284050d",
   760 => x"0402f005",
   761 => x"0d029705",
   762 => x"84808080",
   763 => x"f52d83ff",
   764 => x"f1dc0881",
   765 => x"0583fff1",
   766 => x"dc0c5473",
   767 => x"80d32e09",
   768 => x"8106a338",
   769 => x"800b83ff",
   770 => x"f1dc0c80",
   771 => x"0b83fff1",
   772 => x"cc0c800b",
   773 => x"83fff1e0",
   774 => x"0c800b83",
   775 => x"fff1c80c",
   776 => x"8480809a",
   777 => x"fb0483ff",
   778 => x"f1dc0852",
   779 => x"71812e09",
   780 => x"8106bc38",
   781 => x"83fff1c8",
   782 => x"087481df",
   783 => x"06c90552",
   784 => x"52708025",
   785 => x"8438a711",
   786 => x"5171842b",
   787 => x"71077083",
   788 => x"fff1c80c",
   789 => x"70525283",
   790 => x"72258538",
   791 => x"8a723151",
   792 => x"70108205",
   793 => x"83fff1d4",
   794 => x"0c848080",
   795 => x"9afb0471",
   796 => x"8324a638",
   797 => x"83fff1e0",
   798 => x"087481df",
   799 => x"06c90552",
   800 => x"52708025",
   801 => x"8438a711",
   802 => x"5171842b",
   803 => x"710783ff",
   804 => x"f1e00c84",
   805 => x"80809afb",
   806 => x"0483fff1",
   807 => x"d4088305",
   808 => x"51717124",
   809 => x"a63883ff",
   810 => x"f1cc0874",
   811 => x"81df06c9",
   812 => x"05525270",
   813 => x"80258438",
   814 => x"a7115171",
   815 => x"842b7107",
   816 => x"83fff1cc",
   817 => x"0c848080",
   818 => x"9aba0483",
   819 => x"fff1c808",
   820 => x"ff115253",
   821 => x"70822681",
   822 => x"973883ff",
   823 => x"f1e00810",
   824 => x"81055171",
   825 => x"712480df",
   826 => x"3883fff1",
   827 => x"d8087481",
   828 => x"df06c905",
   829 => x"52527080",
   830 => x"258438a7",
   831 => x"11517184",
   832 => x"2b710770",
   833 => x"83fff1d8",
   834 => x"0c83fff1",
   835 => x"d008ff05",
   836 => x"83fff1d0",
   837 => x"0c5283ff",
   838 => x"f1d00880",
   839 => x"2580dc38",
   840 => x"83fff1cc",
   841 => x"08517171",
   842 => x"84808081",
   843 => x"b72d83ff",
   844 => x"f1cc0881",
   845 => x"0583fff1",
   846 => x"cc0c810b",
   847 => x"83fff1d0",
   848 => x"0c848080",
   849 => x"9afb0483",
   850 => x"fff1d008",
   851 => x"ae3883ff",
   852 => x"f1d80884",
   853 => x"2b7083ff",
   854 => x"f1d80c83",
   855 => x"fff1cc08",
   856 => x"52527171",
   857 => x"84808081",
   858 => x"b72d8480",
   859 => x"809afb04",
   860 => x"86732587",
   861 => x"38848080",
   862 => x"80932d02",
   863 => x"90050d04",
   864 => x"02ec050d",
   865 => x"800bfc80",
   866 => x"0c848080",
   867 => x"b2805184",
   868 => x"808085c5",
   869 => x"2d848080",
   870 => x"93902d83",
   871 => x"ffe08008",
   872 => x"802e8286",
   873 => x"38848080",
   874 => x"b2985184",
   875 => x"808085c5",
   876 => x"2d848080",
   877 => x"9ec02d83",
   878 => x"ffe1a052",
   879 => x"848080b2",
   880 => x"b0518480",
   881 => x"80abf62d",
   882 => x"83ffe080",
   883 => x"08802e81",
   884 => x"cd3883ff",
   885 => x"e1a00b84",
   886 => x"8080b2bc",
   887 => x"52548480",
   888 => x"8085c52d",
   889 => x"80557370",
   890 => x"81055584",
   891 => x"808080f5",
   892 => x"2d5372a0",
   893 => x"2e80e638",
   894 => x"72c00c72",
   895 => x"a32e8184",
   896 => x"387280c7",
   897 => x"2e098106",
   898 => x"8d388480",
   899 => x"8080932d",
   900 => x"8480809c",
   901 => x"b804728a",
   902 => x"2e098106",
   903 => x"8d388480",
   904 => x"80808c2d",
   905 => x"8480809c",
   906 => x"b8047280",
   907 => x"cc2e0981",
   908 => x"06863883",
   909 => x"ffe1a054",
   910 => x"7281df06",
   911 => x"f0057081",
   912 => x"ff065153",
   913 => x"b8732789",
   914 => x"38ef1370",
   915 => x"81ff0651",
   916 => x"5374842b",
   917 => x"73075584",
   918 => x"80809be6",
   919 => x"0472a32e",
   920 => x"a3387370",
   921 => x"81055584",
   922 => x"808080f5",
   923 => x"2d5372a0",
   924 => x"2ef038ff",
   925 => x"14755370",
   926 => x"52548480",
   927 => x"80abf62d",
   928 => x"74fc800c",
   929 => x"73708105",
   930 => x"55848080",
   931 => x"80f52d53",
   932 => x"728a2e09",
   933 => x"8106ed38",
   934 => x"8480809b",
   935 => x"e4048480",
   936 => x"80b2d051",
   937 => x"84808085",
   938 => x"c52d8480",
   939 => x"80b2ec51",
   940 => x"84808085",
   941 => x"c52dae51",
   942 => x"84808085",
   943 => x"a12dbd84",
   944 => x"bf55c008",
   945 => x"70892a70",
   946 => x"81065154",
   947 => x"5472802e",
   948 => x"92387381",
   949 => x"ff065184",
   950 => x"808097e1",
   951 => x"2d848080",
   952 => x"9dbe04ff",
   953 => x"155574ff",
   954 => x"2e098106",
   955 => x"d5388480",
   956 => x"809db604",
   957 => x"02e8050d",
   958 => x"77797b58",
   959 => x"55558053",
   960 => x"727625af",
   961 => x"38747081",
   962 => x"05568480",
   963 => x"8080f52d",
   964 => x"74708105",
   965 => x"56848080",
   966 => x"80f52d52",
   967 => x"5271712e",
   968 => x"89388151",
   969 => x"8480809e",
   970 => x"b5048113",
   971 => x"53848080",
   972 => x"9e800480",
   973 => x"517083ff",
   974 => x"e0800c02",
   975 => x"98050d04",
   976 => x"02d8050d",
   977 => x"800b83ff",
   978 => x"f6940c84",
   979 => x"8080b380",
   980 => x"51848080",
   981 => x"85c52d83",
   982 => x"fff1f052",
   983 => x"80518480",
   984 => x"8095d92d",
   985 => x"83ffe080",
   986 => x"085483ff",
   987 => x"e0800895",
   988 => x"38848080",
   989 => x"b3905184",
   990 => x"808085c5",
   991 => x"2d735584",
   992 => x"8080a6ef",
   993 => x"04848080",
   994 => x"b3a45184",
   995 => x"808085c5",
   996 => x"2d805681",
   997 => x"0b83fff1",
   998 => x"e40c8853",
   999 => x"848080b3",
  1000 => x"bc5283ff",
  1001 => x"f2a65184",
  1002 => x"80809df4",
  1003 => x"2d83ffe0",
  1004 => x"8008762e",
  1005 => x"0981068b",
  1006 => x"3883ffe0",
  1007 => x"800883ff",
  1008 => x"f1e40c88",
  1009 => x"53848080",
  1010 => x"b3c85283",
  1011 => x"fff2c251",
  1012 => x"8480809d",
  1013 => x"f42d83ff",
  1014 => x"e080088b",
  1015 => x"3883ffe0",
  1016 => x"800883ff",
  1017 => x"f1e40c83",
  1018 => x"fff1e408",
  1019 => x"52848080",
  1020 => x"b3d45184",
  1021 => x"808082e3",
  1022 => x"2d83fff1",
  1023 => x"e408802e",
  1024 => x"81cb3883",
  1025 => x"fff5b60b",
  1026 => x"84808080",
  1027 => x"f52d83ff",
  1028 => x"f5b70b84",
  1029 => x"808080f5",
  1030 => x"2d71982b",
  1031 => x"71902b07",
  1032 => x"83fff5b8",
  1033 => x"0b848080",
  1034 => x"80f52d70",
  1035 => x"882b7207",
  1036 => x"83fff5b9",
  1037 => x"0b848080",
  1038 => x"80f52d71",
  1039 => x"0783fff5",
  1040 => x"ee0b8480",
  1041 => x"8080f52d",
  1042 => x"83fff5ef",
  1043 => x"0b848080",
  1044 => x"80f52d71",
  1045 => x"882b0753",
  1046 => x"5f54525a",
  1047 => x"56575573",
  1048 => x"81abaa2e",
  1049 => x"09810695",
  1050 => x"38755184",
  1051 => x"808096db",
  1052 => x"2d83ffe0",
  1053 => x"80085684",
  1054 => x"8080a196",
  1055 => x"047382d4",
  1056 => x"d52e9338",
  1057 => x"848080b3",
  1058 => x"e8518480",
  1059 => x"8085c52d",
  1060 => x"848080a3",
  1061 => x"a2047552",
  1062 => x"848080b4",
  1063 => x"88518480",
  1064 => x"8082e32d",
  1065 => x"83fff1f0",
  1066 => x"52755184",
  1067 => x"808095d9",
  1068 => x"2d83ffe0",
  1069 => x"80085583",
  1070 => x"ffe08008",
  1071 => x"802e85af",
  1072 => x"38848080",
  1073 => x"b4a05184",
  1074 => x"808085c5",
  1075 => x"2d848080",
  1076 => x"b4c85184",
  1077 => x"808082e3",
  1078 => x"2d885384",
  1079 => x"8080b3c8",
  1080 => x"5283fff2",
  1081 => x"c2518480",
  1082 => x"809df42d",
  1083 => x"83ffe080",
  1084 => x"088e3881",
  1085 => x"0b83fff6",
  1086 => x"940c8480",
  1087 => x"80a2ae04",
  1088 => x"88538480",
  1089 => x"80b3bc52",
  1090 => x"83fff2a6",
  1091 => x"51848080",
  1092 => x"9df42d83",
  1093 => x"ffe08008",
  1094 => x"802e9338",
  1095 => x"848080b4",
  1096 => x"e0518480",
  1097 => x"8082e32d",
  1098 => x"848080a3",
  1099 => x"a20483ff",
  1100 => x"f5ee0b84",
  1101 => x"808080f5",
  1102 => x"2d547380",
  1103 => x"d52e0981",
  1104 => x"0680df38",
  1105 => x"83fff5ef",
  1106 => x"0b848080",
  1107 => x"80f52d54",
  1108 => x"7381aa2e",
  1109 => x"09810680",
  1110 => x"c938800b",
  1111 => x"83fff1f0",
  1112 => x"0b848080",
  1113 => x"80f52d56",
  1114 => x"547481e9",
  1115 => x"2e833881",
  1116 => x"547481eb",
  1117 => x"2e8c3880",
  1118 => x"5573752e",
  1119 => x"09810683",
  1120 => x"ee3883ff",
  1121 => x"f1fb0b84",
  1122 => x"808080f5",
  1123 => x"2d597892",
  1124 => x"3883fff1",
  1125 => x"fc0b8480",
  1126 => x"8080f52d",
  1127 => x"5473822e",
  1128 => x"89388055",
  1129 => x"848080a6",
  1130 => x"ef0483ff",
  1131 => x"f1fd0b84",
  1132 => x"808080f5",
  1133 => x"2d7083ff",
  1134 => x"f69c0cff",
  1135 => x"117083ff",
  1136 => x"f6900c54",
  1137 => x"52848080",
  1138 => x"b5805184",
  1139 => x"808082e3",
  1140 => x"2d83fff1",
  1141 => x"fe0b8480",
  1142 => x"8080f52d",
  1143 => x"83fff1ff",
  1144 => x"0b848080",
  1145 => x"80f52d56",
  1146 => x"76057582",
  1147 => x"80290570",
  1148 => x"83fff684",
  1149 => x"0c83fff2",
  1150 => x"800b8480",
  1151 => x"8080f52d",
  1152 => x"7083fff6",
  1153 => x"800c83ff",
  1154 => x"f6940859",
  1155 => x"57587680",
  1156 => x"2e81ec38",
  1157 => x"88538480",
  1158 => x"80b3c852",
  1159 => x"83fff2c2",
  1160 => x"51848080",
  1161 => x"9df42d78",
  1162 => x"5583ffe0",
  1163 => x"800882bf",
  1164 => x"3883fff6",
  1165 => x"9c087084",
  1166 => x"2b83fff5",
  1167 => x"f00c7083",
  1168 => x"fff6980c",
  1169 => x"83fff295",
  1170 => x"0b848080",
  1171 => x"80f52d83",
  1172 => x"fff2940b",
  1173 => x"84808080",
  1174 => x"f52d7182",
  1175 => x"80290583",
  1176 => x"fff2960b",
  1177 => x"84808080",
  1178 => x"f52d7084",
  1179 => x"80802912",
  1180 => x"83fff297",
  1181 => x"0b848080",
  1182 => x"80f52d70",
  1183 => x"81800a29",
  1184 => x"127083ff",
  1185 => x"f1e80c83",
  1186 => x"fff68008",
  1187 => x"712983ff",
  1188 => x"f6840805",
  1189 => x"7083fff6",
  1190 => x"a40c83ff",
  1191 => x"f29d0b84",
  1192 => x"808080f5",
  1193 => x"2d83fff2",
  1194 => x"9c0b8480",
  1195 => x"8080f52d",
  1196 => x"71828029",
  1197 => x"0583fff2",
  1198 => x"9e0b8480",
  1199 => x"8080f52d",
  1200 => x"70848080",
  1201 => x"291283ff",
  1202 => x"f29f0b84",
  1203 => x"808080f5",
  1204 => x"2d70982b",
  1205 => x"81f00a06",
  1206 => x"72057083",
  1207 => x"fff1ec0c",
  1208 => x"fe117e29",
  1209 => x"770583ff",
  1210 => x"f68c0c52",
  1211 => x"5752575d",
  1212 => x"5751525f",
  1213 => x"525c5757",
  1214 => x"57848080",
  1215 => x"a6ed0483",
  1216 => x"fff2820b",
  1217 => x"84808080",
  1218 => x"f52d83ff",
  1219 => x"f2810b84",
  1220 => x"808080f5",
  1221 => x"2d718280",
  1222 => x"29057083",
  1223 => x"fff5f00c",
  1224 => x"70a02983",
  1225 => x"ff057089",
  1226 => x"2a7083ff",
  1227 => x"f6980c83",
  1228 => x"fff2870b",
  1229 => x"84808080",
  1230 => x"f52d83ff",
  1231 => x"f2860b84",
  1232 => x"808080f5",
  1233 => x"2d718280",
  1234 => x"29057083",
  1235 => x"fff1e80c",
  1236 => x"7b71291e",
  1237 => x"7083fff6",
  1238 => x"8c0c7d83",
  1239 => x"fff1ec0c",
  1240 => x"730583ff",
  1241 => x"f6a40c55",
  1242 => x"5e515155",
  1243 => x"55815574",
  1244 => x"83ffe080",
  1245 => x"0c02a805",
  1246 => x"0d0402ec",
  1247 => x"050d7670",
  1248 => x"872c7180",
  1249 => x"ff065556",
  1250 => x"5483fff6",
  1251 => x"94088a38",
  1252 => x"73882c74",
  1253 => x"81ff0654",
  1254 => x"5583fff1",
  1255 => x"f05283ff",
  1256 => x"f6840815",
  1257 => x"51848080",
  1258 => x"95d92d83",
  1259 => x"ffe08008",
  1260 => x"5483ffe0",
  1261 => x"8008802e",
  1262 => x"80c93883",
  1263 => x"fff69408",
  1264 => x"802ea238",
  1265 => x"72842983",
  1266 => x"fff1f005",
  1267 => x"70085253",
  1268 => x"84808096",
  1269 => x"db2d83ff",
  1270 => x"e08008f0",
  1271 => x"0a065384",
  1272 => x"8080a881",
  1273 => x"04721083",
  1274 => x"fff1f005",
  1275 => x"70848080",
  1276 => x"80e02d52",
  1277 => x"53848080",
  1278 => x"97872d83",
  1279 => x"ffe08008",
  1280 => x"53725473",
  1281 => x"83ffe080",
  1282 => x"0c029405",
  1283 => x"0d0402c8",
  1284 => x"050d7f61",
  1285 => x"5f5b800b",
  1286 => x"83fff1ec",
  1287 => x"0883fff6",
  1288 => x"8c08595d",
  1289 => x"5683fff6",
  1290 => x"9408762e",
  1291 => x"8f3883ff",
  1292 => x"f69c0884",
  1293 => x"2b588480",
  1294 => x"80a8c404",
  1295 => x"83fff698",
  1296 => x"08842b58",
  1297 => x"80597878",
  1298 => x"2781dc38",
  1299 => x"788f06a0",
  1300 => x"17575473",
  1301 => x"963883ff",
  1302 => x"f1f05276",
  1303 => x"51811757",
  1304 => x"84808095",
  1305 => x"d92d83ff",
  1306 => x"f1f05680",
  1307 => x"76848080",
  1308 => x"80f52d56",
  1309 => x"5474742e",
  1310 => x"83388154",
  1311 => x"7481e52e",
  1312 => x"819c3881",
  1313 => x"70750655",
  1314 => x"5d73802e",
  1315 => x"8190388b",
  1316 => x"16848080",
  1317 => x"80f52d98",
  1318 => x"065a7981",
  1319 => x"81388b53",
  1320 => x"7d527551",
  1321 => x"8480809d",
  1322 => x"f42d83ff",
  1323 => x"e0800880",
  1324 => x"ed389c16",
  1325 => x"08518480",
  1326 => x"8096db2d",
  1327 => x"83ffe080",
  1328 => x"08841c0c",
  1329 => x"9a168480",
  1330 => x"8080e02d",
  1331 => x"51848080",
  1332 => x"97872d83",
  1333 => x"ffe08008",
  1334 => x"83ffe080",
  1335 => x"08881d0c",
  1336 => x"83ffe080",
  1337 => x"08555583",
  1338 => x"fff69408",
  1339 => x"802ea038",
  1340 => x"94168480",
  1341 => x"8080e02d",
  1342 => x"51848080",
  1343 => x"97872d83",
  1344 => x"ffe08008",
  1345 => x"902b83ff",
  1346 => x"f00a0670",
  1347 => x"16515473",
  1348 => x"881c0c79",
  1349 => x"7b0c7c54",
  1350 => x"848080aa",
  1351 => x"ef048119",
  1352 => x"59848080",
  1353 => x"a8c60483",
  1354 => x"fff69408",
  1355 => x"802ebe38",
  1356 => x"7b518480",
  1357 => x"80a6fa2d",
  1358 => x"83ffe080",
  1359 => x"0883ffe0",
  1360 => x"800880ff",
  1361 => x"fffff806",
  1362 => x"555c7380",
  1363 => x"fffffff8",
  1364 => x"2e9b3883",
  1365 => x"ffe08008",
  1366 => x"fe0583ff",
  1367 => x"f69c0829",
  1368 => x"83fff6a4",
  1369 => x"08055784",
  1370 => x"8080a8c4",
  1371 => x"04805473",
  1372 => x"83ffe080",
  1373 => x"0c02b805",
  1374 => x"0d0402f4",
  1375 => x"050d7470",
  1376 => x"08810571",
  1377 => x"0c700883",
  1378 => x"fff69008",
  1379 => x"06535371",
  1380 => x"93388813",
  1381 => x"08518480",
  1382 => x"80a6fa2d",
  1383 => x"83ffe080",
  1384 => x"0888140c",
  1385 => x"810b83ff",
  1386 => x"e0800c02",
  1387 => x"8c050d04",
  1388 => x"02f0050d",
  1389 => x"75881108",
  1390 => x"fe0583ff",
  1391 => x"f69c0829",
  1392 => x"83fff6a4",
  1393 => x"08117208",
  1394 => x"83fff690",
  1395 => x"08060579",
  1396 => x"55535454",
  1397 => x"84808095",
  1398 => x"d92d83ff",
  1399 => x"e0800853",
  1400 => x"83ffe080",
  1401 => x"08802e83",
  1402 => x"38815372",
  1403 => x"83ffe080",
  1404 => x"0c029005",
  1405 => x"0d0402ec",
  1406 => x"050d7678",
  1407 => x"715483ff",
  1408 => x"f5f45354",
  1409 => x"55848080",
  1410 => x"a88e2d83",
  1411 => x"ffe08008",
  1412 => x"5483ffe0",
  1413 => x"8008802e",
  1414 => x"80ce3884",
  1415 => x"8080b5a4",
  1416 => x"51848080",
  1417 => x"85c52d83",
  1418 => x"fff5f808",
  1419 => x"83ff0589",
  1420 => x"2a558054",
  1421 => x"73752580",
  1422 => x"d1387252",
  1423 => x"83fff5f4",
  1424 => x"51848080",
  1425 => x"abb02d83",
  1426 => x"ffe08008",
  1427 => x"802eaf38",
  1428 => x"83fff5f4",
  1429 => x"51848080",
  1430 => x"aafa2d84",
  1431 => x"80138115",
  1432 => x"55538480",
  1433 => x"80acb404",
  1434 => x"74528480",
  1435 => x"80b5c051",
  1436 => x"84808082",
  1437 => x"e32d7353",
  1438 => x"848080ad",
  1439 => x"8c0483ff",
  1440 => x"e0800853",
  1441 => x"848080ad",
  1442 => x"8c048153",
  1443 => x"7283ffe0",
  1444 => x"800c0294",
  1445 => x"050d0400",
  1446 => x"00ffffff",
  1447 => x"ff00ffff",
  1448 => x"ffff00ff",
  1449 => x"ffffff00",
  1450 => x"53442043",
  1451 => x"4d442025",
  1452 => x"78200000",
  1453 => x"4c424120",
  1454 => x"25782c20",
  1455 => x"00000000",
  1456 => x"27435243",
  1457 => x"27202578",
  1458 => x"20202d3e",
  1459 => x"20000000",
  1460 => x"25780a00",
  1461 => x"434d4435",
  1462 => x"35202564",
  1463 => x"0a000000",
  1464 => x"434d4400",
  1465 => x"696e6974",
  1466 => x"2025640a",
  1467 => x"20200000",
  1468 => x"636d645f",
  1469 => x"434d4438",
  1470 => x"20726573",
  1471 => x"706f6e73",
  1472 => x"653a2025",
  1473 => x"640a0000",
  1474 => x"434d4438",
  1475 => x"5f342072",
  1476 => x"6573706f",
  1477 => x"6e73653a",
  1478 => x"2025640a",
  1479 => x"00000000",
  1480 => x"434d4438",
  1481 => x"202d3e20",
  1482 => x"4e6f7420",
  1483 => x"61205632",
  1484 => x"20636172",
  1485 => x"640a0000",
  1486 => x"5965730a",
  1487 => x"00000000",
  1488 => x"53444843",
  1489 => x"20496e69",
  1490 => x"7469616c",
  1491 => x"697a6174",
  1492 => x"696f6e20",
  1493 => x"6572726f",
  1494 => x"72210a00",
  1495 => x"56322063",
  1496 => x"61726420",
  1497 => x"2d206973",
  1498 => x"20697420",
  1499 => x"53484443",
  1500 => x"3f202000",
  1501 => x"434d4435",
  1502 => x"38202564",
  1503 => x"0a202000",
  1504 => x"434d4435",
  1505 => x"385f3220",
  1506 => x"25640a20",
  1507 => x"20000000",
  1508 => x"4e6f0a00",
  1509 => x"57726974",
  1510 => x"65206661",
  1511 => x"696c6564",
  1512 => x"0a000000",
  1513 => x"434d4439",
  1514 => x"20726573",
  1515 => x"706f6e73",
  1516 => x"653a2025",
  1517 => x"780a0000",
  1518 => x"635f7369",
  1519 => x"7a655f6d",
  1520 => x"756c743a",
  1521 => x"2025642c",
  1522 => x"20726561",
  1523 => x"645f626c",
  1524 => x"5f6c656e",
  1525 => x"3a202564",
  1526 => x"2c206373",
  1527 => x"697a653a",
  1528 => x"2025640a",
  1529 => x"00000000",
  1530 => x"4d756c74",
  1531 => x"2025640a",
  1532 => x"00000000",
  1533 => x"25642062",
  1534 => x"6c6f636b",
  1535 => x"73206f66",
  1536 => x"2073697a",
  1537 => x"65202564",
  1538 => x"0a000000",
  1539 => x"25642062",
  1540 => x"6c6f636b",
  1541 => x"73206f66",
  1542 => x"20353132",
  1543 => x"20627974",
  1544 => x"65730a00",
  1545 => x"53504900",
  1546 => x"41637469",
  1547 => x"76617469",
  1548 => x"6e672043",
  1549 => x"530a0000",
  1550 => x"53656e74",
  1551 => x"20726573",
  1552 => x"65742063",
  1553 => x"6f6d6d61",
  1554 => x"6e640a00",
  1555 => x"43617264",
  1556 => x"20726573",
  1557 => x"706f6e64",
  1558 => x"65642074",
  1559 => x"6f207265",
  1560 => x"7365740a",
  1561 => x"00000000",
  1562 => x"53444843",
  1563 => x"20636172",
  1564 => x"64206465",
  1565 => x"74656374",
  1566 => x"65640a00",
  1567 => x"49455252",
  1568 => x"00000000",
  1569 => x"53442063",
  1570 => x"61726420",
  1571 => x"696e6974",
  1572 => x"69616c69",
  1573 => x"7a617469",
  1574 => x"6f6e2065",
  1575 => x"72726f72",
  1576 => x"210a0000",
  1577 => x"53656e64",
  1578 => x"696e6720",
  1579 => x"636d6431",
  1580 => x"36202862",
  1581 => x"6c6f636b",
  1582 => x"73697a65",
  1583 => x"290a0000",
  1584 => x"53442063",
  1585 => x"61726420",
  1586 => x"73697a65",
  1587 => x"20697320",
  1588 => x"25640a00",
  1589 => x"496e6974",
  1590 => x"20646f6e",
  1591 => x"650a0000",
  1592 => x"52656164",
  1593 => x"20636f6d",
  1594 => x"6d616e64",
  1595 => x"20666169",
  1596 => x"6c656420",
  1597 => x"61742025",
  1598 => x"64202825",
  1599 => x"64290a00",
  1600 => x"496e6974",
  1601 => x"69616c69",
  1602 => x"7a696e67",
  1603 => x"20534420",
  1604 => x"63617264",
  1605 => x"0a000000",
  1606 => x"48756e74",
  1607 => x"696e6720",
  1608 => x"666f7220",
  1609 => x"70617274",
  1610 => x"6974696f",
  1611 => x"6e0a0000",
  1612 => x"4d414e49",
  1613 => x"46455354",
  1614 => x"4d535400",
  1615 => x"50617273",
  1616 => x"696e6720",
  1617 => x"6d616e69",
  1618 => x"66657374",
  1619 => x"0a000000",
  1620 => x"4c6f6164",
  1621 => x"696e6720",
  1622 => x"6d616e69",
  1623 => x"66657374",
  1624 => x"20666169",
  1625 => x"6c65640a",
  1626 => x"00000000",
  1627 => x"426f6f74",
  1628 => x"696e6720",
  1629 => x"66726f6d",
  1630 => x"20525332",
  1631 => x"33322e00",
  1632 => x"52656164",
  1633 => x"696e6720",
  1634 => x"4d42520a",
  1635 => x"00000000",
  1636 => x"52656164",
  1637 => x"206f6620",
  1638 => x"4d425220",
  1639 => x"6661696c",
  1640 => x"65640a00",
  1641 => x"4d425220",
  1642 => x"73756363",
  1643 => x"65737366",
  1644 => x"756c6c79",
  1645 => x"20726561",
  1646 => x"640a0000",
  1647 => x"46415431",
  1648 => x"36202020",
  1649 => x"00000000",
  1650 => x"46415433",
  1651 => x"32202020",
  1652 => x"00000000",
  1653 => x"50617274",
  1654 => x"6974696f",
  1655 => x"6e636f75",
  1656 => x"6e742025",
  1657 => x"640a0000",
  1658 => x"4e6f2070",
  1659 => x"61727469",
  1660 => x"74696f6e",
  1661 => x"20736967",
  1662 => x"6e617475",
  1663 => x"72652066",
  1664 => x"6f756e64",
  1665 => x"0a000000",
  1666 => x"52656164",
  1667 => x"696e6720",
  1668 => x"626f6f74",
  1669 => x"20736563",
  1670 => x"746f7220",
  1671 => x"25640a00",
  1672 => x"52656164",
  1673 => x"20626f6f",
  1674 => x"74207365",
  1675 => x"63746f72",
  1676 => x"2066726f",
  1677 => x"6d206669",
  1678 => x"72737420",
  1679 => x"70617274",
  1680 => x"6974696f",
  1681 => x"6e0a0000",
  1682 => x"48756e74",
  1683 => x"696e6720",
  1684 => x"666f7220",
  1685 => x"66696c65",
  1686 => x"73797374",
  1687 => x"656d0a00",
  1688 => x"556e7375",
  1689 => x"70706f72",
  1690 => x"74656420",
  1691 => x"70617274",
  1692 => x"6974696f",
  1693 => x"6e207479",
  1694 => x"7065210d",
  1695 => x"00000000",
  1696 => x"436c7573",
  1697 => x"74657220",
  1698 => x"73697a65",
  1699 => x"3a202564",
  1700 => x"2c20436c",
  1701 => x"75737465",
  1702 => x"72206d61",
  1703 => x"736b2c20",
  1704 => x"25640a00",
  1705 => x"4f70656e",
  1706 => x"65642066",
  1707 => x"696c652c",
  1708 => x"206c6f61",
  1709 => x"64696e67",
  1710 => x"2e2e2e0a",
  1711 => x"00000000",
  1712 => x"43616e27",
  1713 => x"74206f70",
  1714 => x"656e2025",
  1715 => x"730a0000",
	others => x"00000000"
);

begin

process (clk)
begin
	if (clk'event and clk = '1') then
		if (from_zpu.memAWriteEnable = '1') and (from_zpu.memBWriteEnable = '1') and (from_zpu.memAAddr=from_zpu.memBAddr) and (from_zpu.memAWrite/=from_zpu.memBWrite) then
			report "write collision" severity failure;
		end if;
	
		if (from_zpu.memAWriteEnable = '1') then
			ram(to_integer(unsigned(from_zpu.memAAddr(maxAddrBitBRAM downto 2)))) := from_zpu.memAWrite;
			to_zpu.memARead <= from_zpu.memAWrite;
		else
			to_zpu.memARead <= ram(to_integer(unsigned(from_zpu.memAAddr(maxAddrBitBRAM downto 2))));
		end if;
	end if;
end process;

process (clk)
begin
	if (clk'event and clk = '1') then
		if (from_zpu.memBWriteEnable = '1') then
			ram(to_integer(unsigned(from_zpu.memBAddr(maxAddrBitBRAM downto 2)))) := from_zpu.memBWrite;
			to_zpu.memBRead <= from_zpu.memBWrite;
		else
			to_zpu.memBRead <= ram(to_integer(unsigned(from_zpu.memBAddr(maxAddrBitBRAM downto 2))));
		end if;
	end if;
end process;


end arch;

