-- ZPU
--
-- Copyright 2004-2008 oharboe - �yvind Harboe - oyvind.harboe@zylin.com
-- Modified by Alastair M. Robinson for the ZPUFlex project.
--
-- The FreeBSD license
-- 
-- Redistribution and use in source and binary forms, with or without
-- modification, are permitted provided that the following conditions
-- are met:
-- 
-- 1. Redistributions of source code must retain the above copyright
--    notice, this list of conditions and the following disclaimer.
-- 2. Redistributions in binary form must reproduce the above
--    copyright notice, this list of conditions and the following
--    disclaimer in the documentation and/or other materials
--    provided with the distribution.
-- 
-- THIS SOFTWARE IS PROVIDED BY THE ZPU PROJECT ``AS IS'' AND ANY
-- EXPRESS OR IMPLIED WARRANTIES, INCLUDING, BUT NOT LIMITED TO,
-- THE IMPLIED WARRANTIES OF MERCHANTABILITY AND FITNESS FOR A
-- PARTICULAR PURPOSE ARE DISCLAIMED. IN NO EVENT SHALL THE
-- ZPU PROJECT OR CONTRIBUTORS BE LIABLE FOR ANY DIRECT,
-- INDIRECT, INCIDENTAL, SPECIAL, EXEMPLARY, OR CONSEQUENTIAL DAMAGES
-- (INCLUDING, BUT NOT LIMITED TO, PROCUREMENT OF SUBSTITUTE GOODS
-- OR SERVICES; LOSS OF USE, DATA, OR PROFITS; OR BUSINESS INTERRUPTION)
-- HOWEVER CAUSED AND ON ANY THEORY OF LIABILITY, WHETHER IN CONTRACT,
-- STRICT LIABILITY, OR TORT (INCLUDING NEGLIGENCE OR OTHERWISE)
-- ARISING IN ANY WAY OUT OF THE USE OF THIS SOFTWARE, EVEN IF
-- ADVISED OF THE POSSIBILITY OF SUCH DAMAGE.
-- 
-- The views and conclusions contained in the software and documentation
-- are those of the authors and should not be interpreted as representing
-- official policies, either expressed or implied, of the ZPU Project.

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;


library work;
use work.zpupkg.all;

entity Interrupt_ROM is
generic
	(
		maxAddrBitBRAM : integer := maxAddrBitBRAMLimit -- Specify your actual ROM size to save LEs and unnecessary block RAM usage.
	);
port (
	clk : in std_logic;
	areset : in std_logic := '0';
	from_zpu : in ZPU_ToROM;
	to_zpu : out ZPU_FromROM
);
end Interrupt_ROM;

architecture arch of Interrupt_ROM is

type ram_type is array(natural range 0 to ((2**(maxAddrBitBRAM+1))/4)-1) of std_logic_vector(wordSize-1 downto 0);

shared variable ram : ram_type :=
(
     0 => x"0b0b0b88",
     1 => x"e5040000",
     2 => x"00000000",
     3 => x"00000000",
     4 => x"00000000",
     5 => x"00000000",
     6 => x"00000000",
     7 => x"00000000",
     8 => x"88088c08",
     9 => x"90080b0b",
    10 => x"0b88e108",
    11 => x"2d900c8c",
    12 => x"0c880c04",
    13 => x"00000000",
    14 => x"00000000",
    15 => x"00000000",
    16 => x"71fd0608",
    17 => x"72830609",
    18 => x"81058205",
    19 => x"832b2a83",
    20 => x"ffff0652",
    21 => x"04000000",
    22 => x"00000000",
    23 => x"00000000",
    24 => x"71fd0608",
    25 => x"83ffff73",
    26 => x"83060981",
    27 => x"05820583",
    28 => x"2b2b0906",
    29 => x"7383ffff",
    30 => x"0b0b0b0b",
    31 => x"83a50400",
    32 => x"72098105",
    33 => x"72057373",
    34 => x"09060906",
    35 => x"73097306",
    36 => x"070a8106",
    37 => x"53510400",
    38 => x"00000000",
    39 => x"00000000",
    40 => x"72722473",
    41 => x"732e0753",
    42 => x"51040000",
    43 => x"00000000",
    44 => x"00000000",
    45 => x"00000000",
    46 => x"00000000",
    47 => x"00000000",
    48 => x"71737109",
    49 => x"71068106",
    50 => x"09810572",
    51 => x"0a100a72",
    52 => x"0a100a31",
    53 => x"050a8106",
    54 => x"51515351",
    55 => x"04000000",
    56 => x"72722673",
    57 => x"732e0753",
    58 => x"51040000",
    59 => x"00000000",
    60 => x"00000000",
    61 => x"00000000",
    62 => x"00000000",
    63 => x"00000000",
    64 => x"00000000",
    65 => x"00000000",
    66 => x"00000000",
    67 => x"00000000",
    68 => x"00000000",
    69 => x"00000000",
    70 => x"00000000",
    71 => x"00000000",
    72 => x"0b0b0b88",
    73 => x"ba040000",
    74 => x"00000000",
    75 => x"00000000",
    76 => x"00000000",
    77 => x"00000000",
    78 => x"00000000",
    79 => x"00000000",
    80 => x"720a722b",
    81 => x"0a535104",
    82 => x"00000000",
    83 => x"00000000",
    84 => x"00000000",
    85 => x"00000000",
    86 => x"00000000",
    87 => x"00000000",
    88 => x"72729f06",
    89 => x"0981050b",
    90 => x"0b0b889f",
    91 => x"05040000",
    92 => x"00000000",
    93 => x"00000000",
    94 => x"00000000",
    95 => x"00000000",
    96 => x"72722aff",
    97 => x"739f062a",
    98 => x"0974090a",
    99 => x"8106ff05",
   100 => x"06075351",
   101 => x"04000000",
   102 => x"00000000",
   103 => x"00000000",
   104 => x"71715351",
   105 => x"04067383",
   106 => x"06098105",
   107 => x"8205832b",
   108 => x"0b2b0772",
   109 => x"fc060c51",
   110 => x"51040000",
   111 => x"00000000",
   112 => x"72098105",
   113 => x"72050970",
   114 => x"81050906",
   115 => x"0a810653",
   116 => x"51040000",
   117 => x"00000000",
   118 => x"00000000",
   119 => x"00000000",
   120 => x"72098105",
   121 => x"72050970",
   122 => x"81050906",
   123 => x"0a098106",
   124 => x"53510400",
   125 => x"00000000",
   126 => x"00000000",
   127 => x"00000000",
   128 => x"71098105",
   129 => x"52040000",
   130 => x"00000000",
   131 => x"00000000",
   132 => x"00000000",
   133 => x"00000000",
   134 => x"00000000",
   135 => x"00000000",
   136 => x"72720981",
   137 => x"05055351",
   138 => x"04000000",
   139 => x"00000000",
   140 => x"00000000",
   141 => x"00000000",
   142 => x"00000000",
   143 => x"00000000",
   144 => x"72097206",
   145 => x"73730906",
   146 => x"07535104",
   147 => x"00000000",
   148 => x"00000000",
   149 => x"00000000",
   150 => x"00000000",
   151 => x"00000000",
   152 => x"71fc0608",
   153 => x"72830609",
   154 => x"81058305",
   155 => x"1010102a",
   156 => x"81ff0652",
   157 => x"04000000",
   158 => x"00000000",
   159 => x"00000000",
   160 => x"71fc0608",
   161 => x"0b0b0b91",
   162 => x"9c738306",
   163 => x"10100508",
   164 => x"060b0b0b",
   165 => x"88a20400",
   166 => x"00000000",
   167 => x"00000000",
   168 => x"88088c08",
   169 => x"90087575",
   170 => x"0b0b0b8d",
   171 => x"9f2d5050",
   172 => x"88085690",
   173 => x"0c8c0c88",
   174 => x"0c510400",
   175 => x"00000000",
   176 => x"88088c08",
   177 => x"90087575",
   178 => x"0b0b0b8e",
   179 => x"d12d5050",
   180 => x"88085690",
   181 => x"0c8c0c88",
   182 => x"0c510400",
   183 => x"00000000",
   184 => x"72097081",
   185 => x"0509060a",
   186 => x"8106ff05",
   187 => x"70547106",
   188 => x"73097274",
   189 => x"05ff0506",
   190 => x"07515151",
   191 => x"04000000",
   192 => x"72097081",
   193 => x"0509060a",
   194 => x"098106ff",
   195 => x"05705471",
   196 => x"06730972",
   197 => x"7405ff05",
   198 => x"06075151",
   199 => x"51040000",
   200 => x"05ff0504",
   201 => x"00000000",
   202 => x"00000000",
   203 => x"00000000",
   204 => x"00000000",
   205 => x"00000000",
   206 => x"00000000",
   207 => x"00000000",
   208 => x"04000000",
   209 => x"00000000",
   210 => x"00000000",
   211 => x"00000000",
   212 => x"00000000",
   213 => x"00000000",
   214 => x"00000000",
   215 => x"00000000",
   216 => x"71810552",
   217 => x"04000000",
   218 => x"00000000",
   219 => x"00000000",
   220 => x"00000000",
   221 => x"00000000",
   222 => x"00000000",
   223 => x"00000000",
   224 => x"00000000",
   225 => x"00000000",
   226 => x"00000000",
   227 => x"00000000",
   228 => x"00000000",
   229 => x"00000000",
   230 => x"00000000",
   231 => x"00000000",
   232 => x"02840572",
   233 => x"10100552",
   234 => x"04000000",
   235 => x"00000000",
   236 => x"00000000",
   237 => x"00000000",
   238 => x"00000000",
   239 => x"00000000",
   240 => x"00000000",
   241 => x"00000000",
   242 => x"00000000",
   243 => x"00000000",
   244 => x"00000000",
   245 => x"00000000",
   246 => x"00000000",
   247 => x"00000000",
   248 => x"717105ff",
   249 => x"05715351",
   250 => x"020d0400",
   251 => x"00000000",
   252 => x"00000000",
   253 => x"00000000",
   254 => x"00000000",
   255 => x"00000000",
   256 => x"10101010",
   257 => x"10101010",
   258 => x"10101010",
   259 => x"10101010",
   260 => x"10101010",
   261 => x"10101010",
   262 => x"10101010",
   263 => x"10101053",
   264 => x"51047381",
   265 => x"ff067383",
   266 => x"06098105",
   267 => x"83051010",
   268 => x"102b0772",
   269 => x"fc060c51",
   270 => x"51047272",
   271 => x"80728106",
   272 => x"ff050972",
   273 => x"06057110",
   274 => x"52720a10",
   275 => x"0a5372ed",
   276 => x"38515153",
   277 => x"51040000",
   278 => x"800488da",
   279 => x"04040000",
   280 => x"00000004",
   281 => x"5d88da0b",
   282 => x"8ce904f9",
   283 => x"3d0d797b",
   284 => x"7d0b0b0b",
   285 => x"929c585a",
   286 => x"57548057",
   287 => x"73772589",
   288 => x"38ad5182",
   289 => x"c23f7330",
   290 => x"54738e38",
   291 => x"b00b0b0b",
   292 => x"0b929c34",
   293 => x"811555a0",
   294 => x"39777436",
   295 => x"91ac0553",
   296 => x"72337570",
   297 => x"81055734",
   298 => x"77743554",
   299 => x"73eb3874",
   300 => x"0b0b0b92",
   301 => x"9c2e9138",
   302 => x"ff155574",
   303 => x"33767081",
   304 => x"05583481",
   305 => x"1757e839",
   306 => x"80763476",
   307 => x"880c893d",
   308 => x"0d04f13d",
   309 => x"0d923d57",
   310 => x"80707870",
   311 => x"84055a08",
   312 => x"72415f5d",
   313 => x"587c7084",
   314 => x"055e085a",
   315 => x"805b7998",
   316 => x"2a7a882b",
   317 => x"5b567586",
   318 => x"38775f81",
   319 => x"c3397d80",
   320 => x"2e819d38",
   321 => x"805e7580",
   322 => x"e42e8a38",
   323 => x"7580f82e",
   324 => x"09810689",
   325 => x"38768418",
   326 => x"71085e58",
   327 => x"547580e4",
   328 => x"2e9e3875",
   329 => x"80e4268a",
   330 => x"387580e3",
   331 => x"2ebf3880",
   332 => x"c6397580",
   333 => x"f32ea538",
   334 => x"7580f82e",
   335 => x"8738b839",
   336 => x"8a538339",
   337 => x"90530b0b",
   338 => x"0b92ec52",
   339 => x"7b51fe9b",
   340 => x"3f88080b",
   341 => x"0b0b92ec",
   342 => x"5a55ab39",
   343 => x"76841871",
   344 => x"0870545b",
   345 => x"585480fe",
   346 => x"3f80559a",
   347 => x"39768418",
   348 => x"71085858",
   349 => x"54b639a5",
   350 => x"5180cc3f",
   351 => x"755180c7",
   352 => x"3f821858",
   353 => x"ae3974ff",
   354 => x"16565480",
   355 => x"7425a438",
   356 => x"78708105",
   357 => x"5a337052",
   358 => x"56ad3f81",
   359 => x"1858e739",
   360 => x"75a52e09",
   361 => x"81068538",
   362 => x"815e8839",
   363 => x"7551983f",
   364 => x"81185881",
   365 => x"1b5b837b",
   366 => x"25feb338",
   367 => x"75fea638",
   368 => x"7e880c91",
   369 => x"3d0d04ff",
   370 => x"3d0d7352",
   371 => x"c0087088",
   372 => x"2a708106",
   373 => x"51515170",
   374 => x"802ef138",
   375 => x"71c00c71",
   376 => x"880c833d",
   377 => x"0d04fb3d",
   378 => x"0d807857",
   379 => x"55757084",
   380 => x"05570853",
   381 => x"80547298",
   382 => x"2a73882b",
   383 => x"54527180",
   384 => x"2ea238c0",
   385 => x"0870882a",
   386 => x"70810651",
   387 => x"51517080",
   388 => x"2ef13871",
   389 => x"c00c8115",
   390 => x"81155555",
   391 => x"837425d6",
   392 => x"3871ca38",
   393 => x"74880c87",
   394 => x"3d0d0471",
   395 => x"88e10c04",
   396 => x"ffb00888",
   397 => x"0c04810b",
   398 => x"ffb00c04",
   399 => x"800bffb0",
   400 => x"0c04ff3d",
   401 => x"0df63fe8",
   402 => x"3f93ac08",
   403 => x"81327093",
   404 => x"ac0c5271",
   405 => x"802e8638",
   406 => x"91c05184",
   407 => x"3991cc51",
   408 => x"ff843fd2",
   409 => x"3f833d0d",
   410 => x"04803d0d",
   411 => x"800b93ac",
   412 => x"0c91d851",
   413 => x"fef03f80",
   414 => x"0bf8840c",
   415 => x"868da00b",
   416 => x"f8880c91",
   417 => x"f051fede",
   418 => x"3f8cc251",
   419 => x"ff9d3fff",
   420 => x"a53f9288",
   421 => x"51fecf3f",
   422 => x"810bf880",
   423 => x"0cff3994",
   424 => x"0802940c",
   425 => x"f93d0d80",
   426 => x"0b9408fc",
   427 => x"050c9408",
   428 => x"88050880",
   429 => x"25ab3894",
   430 => x"08880508",
   431 => x"30940888",
   432 => x"050c800b",
   433 => x"9408f405",
   434 => x"0c9408fc",
   435 => x"05088838",
   436 => x"810b9408",
   437 => x"f4050c94",
   438 => x"08f40508",
   439 => x"9408fc05",
   440 => x"0c94088c",
   441 => x"05088025",
   442 => x"ab389408",
   443 => x"8c050830",
   444 => x"94088c05",
   445 => x"0c800b94",
   446 => x"08f0050c",
   447 => x"9408fc05",
   448 => x"08883881",
   449 => x"0b9408f0",
   450 => x"050c9408",
   451 => x"f0050894",
   452 => x"08fc050c",
   453 => x"80539408",
   454 => x"8c050852",
   455 => x"94088805",
   456 => x"085181a7",
   457 => x"3f880870",
   458 => x"9408f805",
   459 => x"0c549408",
   460 => x"fc050880",
   461 => x"2e8c3894",
   462 => x"08f80508",
   463 => x"309408f8",
   464 => x"050c9408",
   465 => x"f8050870",
   466 => x"880c5489",
   467 => x"3d0d940c",
   468 => x"04940802",
   469 => x"940cfb3d",
   470 => x"0d800b94",
   471 => x"08fc050c",
   472 => x"94088805",
   473 => x"08802593",
   474 => x"38940888",
   475 => x"05083094",
   476 => x"0888050c",
   477 => x"810b9408",
   478 => x"fc050c94",
   479 => x"088c0508",
   480 => x"80258c38",
   481 => x"94088c05",
   482 => x"08309408",
   483 => x"8c050c81",
   484 => x"5394088c",
   485 => x"05085294",
   486 => x"08880508",
   487 => x"51ad3f88",
   488 => x"08709408",
   489 => x"f8050c54",
   490 => x"9408fc05",
   491 => x"08802e8c",
   492 => x"389408f8",
   493 => x"05083094",
   494 => x"08f8050c",
   495 => x"9408f805",
   496 => x"0870880c",
   497 => x"54873d0d",
   498 => x"940c0494",
   499 => x"0802940c",
   500 => x"fd3d0d81",
   501 => x"0b9408fc",
   502 => x"050c800b",
   503 => x"9408f805",
   504 => x"0c94088c",
   505 => x"05089408",
   506 => x"88050827",
   507 => x"ac389408",
   508 => x"fc050880",
   509 => x"2ea33880",
   510 => x"0b94088c",
   511 => x"05082499",
   512 => x"3894088c",
   513 => x"05081094",
   514 => x"088c050c",
   515 => x"9408fc05",
   516 => x"08109408",
   517 => x"fc050cc9",
   518 => x"399408fc",
   519 => x"0508802e",
   520 => x"80c93894",
   521 => x"088c0508",
   522 => x"94088805",
   523 => x"0826a138",
   524 => x"94088805",
   525 => x"0894088c",
   526 => x"05083194",
   527 => x"0888050c",
   528 => x"9408f805",
   529 => x"089408fc",
   530 => x"05080794",
   531 => x"08f8050c",
   532 => x"9408fc05",
   533 => x"08812a94",
   534 => x"08fc050c",
   535 => x"94088c05",
   536 => x"08812a94",
   537 => x"088c050c",
   538 => x"ffaf3994",
   539 => x"08900508",
   540 => x"802e8f38",
   541 => x"94088805",
   542 => x"08709408",
   543 => x"f4050c51",
   544 => x"8d399408",
   545 => x"f8050870",
   546 => x"9408f405",
   547 => x"0c519408",
   548 => x"f4050888",
   549 => x"0c853d0d",
   550 => x"940c0400",
   551 => x"00ffffff",
   552 => x"ff00ffff",
   553 => x"ffff00ff",
   554 => x"ffffff00",
   555 => x"30313233",
   556 => x"34353637",
   557 => x"38394142",
   558 => x"43444546",
   559 => x"00000000",
   560 => x"5469636b",
   561 => x"2e2e2e0a",
   562 => x"00000000",
   563 => x"546f636b",
   564 => x"2e2e2e0a",
   565 => x"00000000",
   566 => x"53657474",
   567 => x"696e6720",
   568 => x"75702074",
   569 => x"696d6572",
   570 => x"2e2e2e0a",
   571 => x"00000000",
   572 => x"456e6162",
   573 => x"6c696e67",
   574 => x"20696e74",
   575 => x"65727275",
   576 => x"7074732e",
   577 => x"2e2e0a00",
   578 => x"456e6162",
   579 => x"6c696e67",
   580 => x"2074696d",
   581 => x"65722e2e",
   582 => x"2e0a002e",
	others => x"00000000"
);

begin

process (clk)
begin
	if (clk'event and clk = '1') then
		if (from_zpu.memAWriteEnable = '1') and (from_zpu.memBWriteEnable = '1') and (from_zpu.memAAddr=from_zpu.memBAddr) and (from_zpu.memAWrite/=from_zpu.memBWrite) then
			report "write collision" severity failure;
		end if;
	
		if (from_zpu.memAWriteEnable = '1') then
			ram(to_integer(unsigned(from_zpu.memAAddr(maxAddrBitBRAM downto 2)))) := from_zpu.memAWrite;
			to_zpu.memARead <= from_zpu.memAWrite;
		else
			to_zpu.memARead <= ram(to_integer(unsigned(from_zpu.memAAddr(maxAddrBitBRAM downto 2))));
		end if;
	end if;
end process;

process (clk)
begin
	if (clk'event and clk = '1') then
		if (from_zpu.memBWriteEnable = '1') then
			ram(to_integer(unsigned(from_zpu.memBAddr(maxAddrBitBRAM downto 2)))) := from_zpu.memBWrite;
			to_zpu.memBRead <= from_zpu.memBWrite;
		else
			to_zpu.memBRead <= ram(to_integer(unsigned(from_zpu.memBAddr(maxAddrBitBRAM downto 2))));
		end if;
	end if;
end process;


end arch;

