-- ZPU
--
-- Copyright 2004-2008 oharboe - �yvind Harboe - oyvind.harboe@zylin.com
-- Modified by Alastair M. Robinson for the ZPUFlex project.
--
-- The FreeBSD license
-- 
-- Redistribution and use in source and binary forms, with or without
-- modification, are permitted provided that the following conditions
-- are met:
-- 
-- 1. Redistributions of source code must retain the above copyright
--    notice, this list of conditions and the following disclaimer.
-- 2. Redistributions in binary form must reproduce the above
--    copyright notice, this list of conditions and the following
--    disclaimer in the documentation and/or other materials
--    provided with the distribution.
-- 
-- THIS SOFTWARE IS PROVIDED BY THE ZPU PROJECT ``AS IS'' AND ANY
-- EXPRESS OR IMPLIED WARRANTIES, INCLUDING, BUT NOT LIMITED TO,
-- THE IMPLIED WARRANTIES OF MERCHANTABILITY AND FITNESS FOR A
-- PARTICULAR PURPOSE ARE DISCLAIMED. IN NO EVENT SHALL THE
-- ZPU PROJECT OR CONTRIBUTORS BE LIABLE FOR ANY DIRECT,
-- INDIRECT, INCIDENTAL, SPECIAL, EXEMPLARY, OR CONSEQUENTIAL DAMAGES
-- (INCLUDING, BUT NOT LIMITED TO, PROCUREMENT OF SUBSTITUTE GOODS
-- OR SERVICES; LOSS OF USE, DATA, OR PROFITS; OR BUSINESS INTERRUPTION)
-- HOWEVER CAUSED AND ON ANY THEORY OF LIABILITY, WHETHER IN CONTRACT,
-- STRICT LIABILITY, OR TORT (INCLUDING NEGLIGENCE OR OTHERWISE)
-- ARISING IN ANY WAY OUT OF THE USE OF THIS SOFTWARE, EVEN IF
-- ADVISED OF THE POSSIBILITY OF SUCH DAMAGE.
-- 
-- The views and conclusions contained in the software and documentation
-- are those of the authors and should not be interpreted as representing
-- official policies, either expressed or implied, of the ZPU Project.

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;


library work;
use work.zpu_config.all;
use work.zpupkg.all;

entity SDBootstrap_ROM is
generic
	(
		maxAddrBit : integer := maxAddrBitBRAMLimit -- Specify your actual ROM size to save LEs and unnecessary block RAM usage.
	);
port (
	clk : in std_logic;
	areset : in std_logic := '0';
	from_zpu : in ZPU_ToROM;
	to_zpu : out ZPU_FromROM
);
end SDBootstrap_ROM;

architecture arch of SDBootstrap_ROM is

type ram_type is array(natural range 0 to ((2**(maxAddrBit+1))/4)-1) of std_logic_vector(wordSize-1 downto 0);

shared variable ram : ram_type :=
(
     0 => x"0ba08080",
     1 => x"e2040000",
     2 => x"8004a080",
     3 => x"808a0471",
     4 => x"fd060872",
     5 => x"83060981",
     6 => x"05820583",
     7 => x"2b2a83ff",
     8 => x"ff065204",
     9 => x"71fc0608",
    10 => x"72830609",
    11 => x"81058305",
    12 => x"1010102a",
    13 => x"81ff0652",
    14 => x"0471fc06",
    15 => x"080ba080",
    16 => x"97fc7383",
    17 => x"06101005",
    18 => x"08067381",
    19 => x"ff067383",
    20 => x"06098105",
    21 => x"83051010",
    22 => x"102b0772",
    23 => x"fc060c51",
    24 => x"5104a080",
    25 => x"808a0ba0",
    26 => x"8087f704",
    27 => x"0002f405",
    28 => x"0d747671",
    29 => x"81ff06d4",
    30 => x"0c535383",
    31 => x"fff09008",
    32 => x"85387189",
    33 => x"2b527198",
    34 => x"2ad40c71",
    35 => x"902a7081",
    36 => x"ff06d40c",
    37 => x"5171882a",
    38 => x"7081ff06",
    39 => x"d40c5171",
    40 => x"81ff06d4",
    41 => x"0c72902a",
    42 => x"7081ff06",
    43 => x"d40c51d4",
    44 => x"087081ff",
    45 => x"06515182",
    46 => x"b8bf5270",
    47 => x"81ff2e09",
    48 => x"81069438",
    49 => x"81ff0bd4",
    50 => x"0cd40870",
    51 => x"81ff06ff",
    52 => x"14545151",
    53 => x"71e53870",
    54 => x"83ffe080",
    55 => x"0c028c05",
    56 => x"0d0402fc",
    57 => x"050d81c7",
    58 => x"5181ff0b",
    59 => x"d40cff11",
    60 => x"51708025",
    61 => x"f4380284",
    62 => x"050d0402",
    63 => x"f0050da0",
    64 => x"8081e22d",
    65 => x"819c9f53",
    66 => x"805287fc",
    67 => x"80f751a0",
    68 => x"8080ed2d",
    69 => x"83ffe080",
    70 => x"085483ff",
    71 => x"e0800881",
    72 => x"2e098106",
    73 => x"ab3881ff",
    74 => x"0bd40c82",
    75 => x"0a52849c",
    76 => x"80e951a0",
    77 => x"8080ed2d",
    78 => x"83ffe080",
    79 => x"088d3881",
    80 => x"ff0bd40c",
    81 => x"7353a080",
    82 => x"82d704a0",
    83 => x"8081e22d",
    84 => x"ff135372",
    85 => x"ffb23872",
    86 => x"83ffe080",
    87 => x"0c029005",
    88 => x"0d0402f4",
    89 => x"050d81ff",
    90 => x"0bd40c93",
    91 => x"53805287",
    92 => x"fc80c151",
    93 => x"a08080ed",
    94 => x"2d83ffe0",
    95 => x"80088d38",
    96 => x"81ff0bd4",
    97 => x"0c8153a0",
    98 => x"80839704",
    99 => x"a08081e2",
   100 => x"2dff1353",
   101 => x"72d73872",
   102 => x"83ffe080",
   103 => x"0c028c05",
   104 => x"0d0402f0",
   105 => x"050da080",
   106 => x"81e22d83",
   107 => x"aa52849c",
   108 => x"80c851a0",
   109 => x"8080ed2d",
   110 => x"83ffe080",
   111 => x"08812e09",
   112 => x"81069038",
   113 => x"d8087083",
   114 => x"ffff0651",
   115 => x"537283aa",
   116 => x"2e9938a0",
   117 => x"8082e22d",
   118 => x"a08083e4",
   119 => x"048154a0",
   120 => x"8084c504",
   121 => x"8054a080",
   122 => x"84c50481",
   123 => x"ff0bd40c",
   124 => x"b153a080",
   125 => x"81fb2d83",
   126 => x"ffe08008",
   127 => x"802eb738",
   128 => x"805287fc",
   129 => x"80fa51a0",
   130 => x"8080ed2d",
   131 => x"83ffe080",
   132 => x"08a43881",
   133 => x"ff0bd40c",
   134 => x"d408d808",
   135 => x"71862a70",
   136 => x"810683ff",
   137 => x"e0800853",
   138 => x"51525553",
   139 => x"72802e95",
   140 => x"38a08083",
   141 => x"dd047282",
   142 => x"2effa938",
   143 => x"ff135372",
   144 => x"ffb03872",
   145 => x"547383ff",
   146 => x"e0800c02",
   147 => x"90050d04",
   148 => x"02f4050d",
   149 => x"810b83ff",
   150 => x"f0900cd0",
   151 => x"08708f2a",
   152 => x"70810651",
   153 => x"515372f3",
   154 => x"3872d00c",
   155 => x"a08081e2",
   156 => x"2dd00870",
   157 => x"8f2a7081",
   158 => x"06515153",
   159 => x"72f33881",
   160 => x"0bd00c87",
   161 => x"53805284",
   162 => x"d480c051",
   163 => x"a08080ed",
   164 => x"2d83ffe0",
   165 => x"8008812e",
   166 => x"96387282",
   167 => x"2e098106",
   168 => x"88388053",
   169 => x"a08085e7",
   170 => x"04ff1353",
   171 => x"72d738a0",
   172 => x"8083a22d",
   173 => x"83ffe080",
   174 => x"0883fff0",
   175 => x"900c8152",
   176 => x"87fc80d0",
   177 => x"51a08080",
   178 => x"ed2d81ff",
   179 => x"0bd40cd0",
   180 => x"08708f2a",
   181 => x"70810651",
   182 => x"515372f3",
   183 => x"3872d00c",
   184 => x"81ff0bd4",
   185 => x"0c815372",
   186 => x"83ffe080",
   187 => x"0c028c05",
   188 => x"0d04800b",
   189 => x"83ffe080",
   190 => x"0c0402e8",
   191 => x"050d7855",
   192 => x"8056d008",
   193 => x"708f2a70",
   194 => x"81065151",
   195 => x"5372f338",
   196 => x"82810bd0",
   197 => x"0c81ff0b",
   198 => x"d40c7752",
   199 => x"87fc80d1",
   200 => x"51a08080",
   201 => x"ed2d83ff",
   202 => x"e0800880",
   203 => x"d23880db",
   204 => x"c6df5481",
   205 => x"ff0bd40c",
   206 => x"d4087081",
   207 => x"ff065153",
   208 => x"7281fe2e",
   209 => x"0981069b",
   210 => x"3880ff54",
   211 => x"d8087570",
   212 => x"8405570c",
   213 => x"ff145473",
   214 => x"8025f138",
   215 => x"8156a080",
   216 => x"86e904ff",
   217 => x"145473cb",
   218 => x"3881ff0b",
   219 => x"d40cd008",
   220 => x"708f2a70",
   221 => x"81065151",
   222 => x"5372f338",
   223 => x"72d00c75",
   224 => x"83ffe080",
   225 => x"0c029805",
   226 => x"0d0402f4",
   227 => x"050d7470",
   228 => x"882a83fe",
   229 => x"80067072",
   230 => x"982a0772",
   231 => x"882b87fc",
   232 => x"80800673",
   233 => x"982b81f0",
   234 => x"0a067173",
   235 => x"070783ff",
   236 => x"e0800c56",
   237 => x"51535102",
   238 => x"8c050d04",
   239 => x"02f4050d",
   240 => x"029205a0",
   241 => x"80808f2d",
   242 => x"70882a71",
   243 => x"882b0770",
   244 => x"83ffff06",
   245 => x"83ffe080",
   246 => x"0c525202",
   247 => x"8c050d04",
   248 => x"02f8050d",
   249 => x"7370902b",
   250 => x"71902a07",
   251 => x"83ffe080",
   252 => x"0c520288",
   253 => x"050d0402",
   254 => x"ec050d80",
   255 => x"0b870a0c",
   256 => x"a08084d0",
   257 => x"2d83ffe0",
   258 => x"8008802e",
   259 => x"81d138a0",
   260 => x"808ab32d",
   261 => x"83ffe090",
   262 => x"52a08098",
   263 => x"8c51a080",
   264 => x"95b82d83",
   265 => x"ffe08008",
   266 => x"802e81b3",
   267 => x"3883ffe0",
   268 => x"90548055",
   269 => x"73708105",
   270 => x"55a08080",
   271 => x"a42d5372",
   272 => x"a02e80de",
   273 => x"3872a32e",
   274 => x"80fd3872",
   275 => x"80c72e09",
   276 => x"81068b38",
   277 => x"a0808088",
   278 => x"2da08088",
   279 => x"fe04728a",
   280 => x"2e098106",
   281 => x"8b38a080",
   282 => x"808a2da0",
   283 => x"8088fe04",
   284 => x"7280cc2e",
   285 => x"09810686",
   286 => x"3883ffe0",
   287 => x"90547281",
   288 => x"df06f005",
   289 => x"7081ff06",
   290 => x"5153b873",
   291 => x"278938ef",
   292 => x"137081ff",
   293 => x"06515374",
   294 => x"842b7307",
   295 => x"55a08088",
   296 => x"b40472a3",
   297 => x"2ea13873",
   298 => x"70810555",
   299 => x"a08080a4",
   300 => x"2d5372a0",
   301 => x"2ef138ff",
   302 => x"14755370",
   303 => x"5254a080",
   304 => x"95b82d74",
   305 => x"870a0c73",
   306 => x"70810555",
   307 => x"a08080a4",
   308 => x"2d53728a",
   309 => x"2e098106",
   310 => x"ee38a080",
   311 => x"88b20480",
   312 => x"0b83ffe0",
   313 => x"800c0294",
   314 => x"050d0402",
   315 => x"e8050d77",
   316 => x"797b5855",
   317 => x"55805372",
   318 => x"7625ab38",
   319 => x"74708105",
   320 => x"56a08080",
   321 => x"a42d7470",
   322 => x"810556a0",
   323 => x"8080a42d",
   324 => x"52527171",
   325 => x"2e883881",
   326 => x"51a0808a",
   327 => x"a8048113",
   328 => x"53a08089",
   329 => x"f7048051",
   330 => x"7083ffe0",
   331 => x"800c0298",
   332 => x"050d0402",
   333 => x"d8050dff",
   334 => x"0b83fff4",
   335 => x"bc0c800b",
   336 => x"83fff4d0",
   337 => x"0c83fff0",
   338 => x"a8528051",
   339 => x"a08085fa",
   340 => x"2d83ffe0",
   341 => x"80085583",
   342 => x"ffe08008",
   343 => x"802e86d3",
   344 => x"38805681",
   345 => x"0b83fff0",
   346 => x"9c0c8853",
   347 => x"a0809898",
   348 => x"5283fff0",
   349 => x"de51a080",
   350 => x"89eb2d83",
   351 => x"ffe08008",
   352 => x"762e0981",
   353 => x"068b3883",
   354 => x"ffe08008",
   355 => x"83fff09c",
   356 => x"0c8853a0",
   357 => x"8098a452",
   358 => x"83fff0fa",
   359 => x"51a08089",
   360 => x"eb2d83ff",
   361 => x"e080088b",
   362 => x"3883ffe0",
   363 => x"800883ff",
   364 => x"f09c0c83",
   365 => x"fff09c08",
   366 => x"802e819c",
   367 => x"3883fff3",
   368 => x"ee0ba080",
   369 => x"80a42d83",
   370 => x"fff3ef0b",
   371 => x"a08080a4",
   372 => x"2d71982b",
   373 => x"71902b07",
   374 => x"83fff3f0",
   375 => x"0ba08080",
   376 => x"a42d7088",
   377 => x"2b720783",
   378 => x"fff3f10b",
   379 => x"a08080a4",
   380 => x"2d710783",
   381 => x"fff4a60b",
   382 => x"a08080a4",
   383 => x"2d83fff4",
   384 => x"a70ba080",
   385 => x"80a42d71",
   386 => x"882b0753",
   387 => x"5f54525a",
   388 => x"56575573",
   389 => x"81abaa2e",
   390 => x"09810693",
   391 => x"387551a0",
   392 => x"80878a2d",
   393 => x"83ffe080",
   394 => x"0856a080",
   395 => x"8cbc0480",
   396 => x"557382d4",
   397 => x"d52e0981",
   398 => x"0684f838",
   399 => x"83fff0a8",
   400 => x"527551a0",
   401 => x"8085fa2d",
   402 => x"83ffe080",
   403 => x"085583ff",
   404 => x"e0800880",
   405 => x"2e84dc38",
   406 => x"8853a080",
   407 => x"98a45283",
   408 => x"fff0fa51",
   409 => x"a08089eb",
   410 => x"2d83ffe0",
   411 => x"80088d38",
   412 => x"810b83ff",
   413 => x"f4d00ca0",
   414 => x"808d9c04",
   415 => x"8853a080",
   416 => x"98985283",
   417 => x"fff0de51",
   418 => x"a08089eb",
   419 => x"2d805583",
   420 => x"ffe08008",
   421 => x"752e0981",
   422 => x"06849838",
   423 => x"83fff4a6",
   424 => x"0ba08080",
   425 => x"a42d5473",
   426 => x"80d52e09",
   427 => x"810680db",
   428 => x"3883fff4",
   429 => x"a70ba080",
   430 => x"80a42d54",
   431 => x"7381aa2e",
   432 => x"09810680",
   433 => x"c638800b",
   434 => x"83fff0a8",
   435 => x"0ba08080",
   436 => x"a42d5654",
   437 => x"7481e92e",
   438 => x"83388154",
   439 => x"7481eb2e",
   440 => x"8c388055",
   441 => x"73752e09",
   442 => x"810683c7",
   443 => x"3883fff0",
   444 => x"b30ba080",
   445 => x"80a42d55",
   446 => x"74913883",
   447 => x"fff0b40b",
   448 => x"a08080a4",
   449 => x"2d547382",
   450 => x"2e883880",
   451 => x"55a08091",
   452 => x"b30483ff",
   453 => x"f0b50ba0",
   454 => x"8080a42d",
   455 => x"7083fff4",
   456 => x"d80cff05",
   457 => x"83fff4cc",
   458 => x"0c83fff0",
   459 => x"b60ba080",
   460 => x"80a42d83",
   461 => x"fff0b70b",
   462 => x"a08080a4",
   463 => x"2d587605",
   464 => x"77828029",
   465 => x"057083ff",
   466 => x"f4c00c83",
   467 => x"fff0b80b",
   468 => x"a08080a4",
   469 => x"2d7083ff",
   470 => x"f4b80c83",
   471 => x"fff4d008",
   472 => x"59575876",
   473 => x"802e81df",
   474 => x"388853a0",
   475 => x"8098a452",
   476 => x"83fff0fa",
   477 => x"51a08089",
   478 => x"eb2d83ff",
   479 => x"e0800882",
   480 => x"b23883ff",
   481 => x"f4d80870",
   482 => x"842b83ff",
   483 => x"f4a80c70",
   484 => x"83fff4d4",
   485 => x"0c83fff0",
   486 => x"cd0ba080",
   487 => x"80a42d83",
   488 => x"fff0cc0b",
   489 => x"a08080a4",
   490 => x"2d718280",
   491 => x"290583ff",
   492 => x"f0ce0ba0",
   493 => x"8080a42d",
   494 => x"70848080",
   495 => x"291283ff",
   496 => x"f0cf0ba0",
   497 => x"8080a42d",
   498 => x"7081800a",
   499 => x"29127083",
   500 => x"fff0a00c",
   501 => x"83fff4b8",
   502 => x"08712983",
   503 => x"fff4c008",
   504 => x"057083ff",
   505 => x"f4e00c83",
   506 => x"fff0d50b",
   507 => x"a08080a4",
   508 => x"2d83fff0",
   509 => x"d40ba080",
   510 => x"80a42d71",
   511 => x"82802905",
   512 => x"83fff0d6",
   513 => x"0ba08080",
   514 => x"a42d7084",
   515 => x"80802912",
   516 => x"83fff0d7",
   517 => x"0ba08080",
   518 => x"a42d7098",
   519 => x"2b81f00a",
   520 => x"06720570",
   521 => x"83fff0a4",
   522 => x"0cfe117e",
   523 => x"29770583",
   524 => x"fff4c80c",
   525 => x"52595243",
   526 => x"545e5152",
   527 => x"59525d57",
   528 => x"5957a080",
   529 => x"91b10483",
   530 => x"fff0ba0b",
   531 => x"a08080a4",
   532 => x"2d83fff0",
   533 => x"b90ba080",
   534 => x"80a42d71",
   535 => x"82802905",
   536 => x"7083fff4",
   537 => x"a80c70a0",
   538 => x"2983ff05",
   539 => x"70892a70",
   540 => x"83fff4d4",
   541 => x"0c83fff0",
   542 => x"bf0ba080",
   543 => x"80a42d83",
   544 => x"fff0be0b",
   545 => x"a08080a4",
   546 => x"2d718280",
   547 => x"29057083",
   548 => x"fff0a00c",
   549 => x"7b71291e",
   550 => x"7083fff4",
   551 => x"c80c7d83",
   552 => x"fff0a40c",
   553 => x"730583ff",
   554 => x"f4e00c55",
   555 => x"5e515155",
   556 => x"55815574",
   557 => x"83ffe080",
   558 => x"0c02a805",
   559 => x"0d0402ec",
   560 => x"050d7670",
   561 => x"872c7180",
   562 => x"ff065755",
   563 => x"5383fff4",
   564 => x"d0088a38",
   565 => x"72882c73",
   566 => x"81ff0656",
   567 => x"547383ff",
   568 => x"f4bc082e",
   569 => x"a83883ff",
   570 => x"f0a85283",
   571 => x"fff4c008",
   572 => x"1451a080",
   573 => x"85fa2d83",
   574 => x"ffe08008",
   575 => x"5383ffe0",
   576 => x"8008802e",
   577 => x"80cb3873",
   578 => x"83fff4bc",
   579 => x"0c83fff4",
   580 => x"d008802e",
   581 => x"a0387484",
   582 => x"2983fff0",
   583 => x"a8057008",
   584 => x"5253a080",
   585 => x"878a2d83",
   586 => x"ffe08008",
   587 => x"f00a0655",
   588 => x"a08092cf",
   589 => x"04741083",
   590 => x"fff0a805",
   591 => x"70a08080",
   592 => x"8f2d5253",
   593 => x"a08087bc",
   594 => x"2d83ffe0",
   595 => x"80085574",
   596 => x"537283ff",
   597 => x"e0800c02",
   598 => x"94050d04",
   599 => x"02cc050d",
   600 => x"7e605e5b",
   601 => x"8056ff0b",
   602 => x"83fff4bc",
   603 => x"0c83fff0",
   604 => x"a40883ff",
   605 => x"f4c80856",
   606 => x"5a83fff4",
   607 => x"d008762e",
   608 => x"8e3883ff",
   609 => x"f4d80884",
   610 => x"2b58a080",
   611 => x"93970483",
   612 => x"fff4d408",
   613 => x"842b5880",
   614 => x"59787827",
   615 => x"81c93878",
   616 => x"8f06a017",
   617 => x"57547395",
   618 => x"3883fff0",
   619 => x"a8527451",
   620 => x"811555a0",
   621 => x"8085fa2d",
   622 => x"83fff0a8",
   623 => x"568076a0",
   624 => x"8080a42d",
   625 => x"55577377",
   626 => x"2e833881",
   627 => x"577381e5",
   628 => x"2e818c38",
   629 => x"81707806",
   630 => x"555c7380",
   631 => x"2e818038",
   632 => x"8b16a080",
   633 => x"80a42d98",
   634 => x"06577680",
   635 => x"f2388b53",
   636 => x"7c527551",
   637 => x"a08089eb",
   638 => x"2d83ffe0",
   639 => x"800880df",
   640 => x"389c1608",
   641 => x"51a08087",
   642 => x"8a2d83ff",
   643 => x"e0800884",
   644 => x"1c0c9a16",
   645 => x"a080808f",
   646 => x"2d51a080",
   647 => x"87bc2d83",
   648 => x"ffe08008",
   649 => x"83ffe080",
   650 => x"08555583",
   651 => x"fff4d008",
   652 => x"802e9e38",
   653 => x"9416a080",
   654 => x"808f2d51",
   655 => x"a08087bc",
   656 => x"2d83ffe0",
   657 => x"8008902b",
   658 => x"83fff00a",
   659 => x"06701651",
   660 => x"5473881c",
   661 => x"0c767b0c",
   662 => x"7b54a080",
   663 => x"95ad0481",
   664 => x"1959a080",
   665 => x"93990483",
   666 => x"fff4d008",
   667 => x"802ebc38",
   668 => x"7951a080",
   669 => x"91be2d83",
   670 => x"ffe08008",
   671 => x"83ffe080",
   672 => x"0880ffff",
   673 => x"fff80655",
   674 => x"5a7380ff",
   675 => x"fffff82e",
   676 => x"9a3883ff",
   677 => x"e08008fe",
   678 => x"0583fff4",
   679 => x"d8082983",
   680 => x"fff4e008",
   681 => x"0555a080",
   682 => x"93970480",
   683 => x"547383ff",
   684 => x"e0800c02",
   685 => x"b4050d04",
   686 => x"02e4050d",
   687 => x"79795383",
   688 => x"fff4ac52",
   689 => x"55a08092",
   690 => x"dc2d83ff",
   691 => x"e0800881",
   692 => x"ff067055",
   693 => x"5372802e",
   694 => x"81853883",
   695 => x"fff4b008",
   696 => x"83ff0589",
   697 => x"2a578070",
   698 => x"55567577",
   699 => x"2580ee38",
   700 => x"83fff4b4",
   701 => x"08fe0583",
   702 => x"fff4d808",
   703 => x"2983fff4",
   704 => x"e0081175",
   705 => x"83fff4cc",
   706 => x"08060576",
   707 => x"545253a0",
   708 => x"8085fa2d",
   709 => x"83ffe080",
   710 => x"08802eb6",
   711 => x"38811470",
   712 => x"83fff4cc",
   713 => x"08065454",
   714 => x"72963883",
   715 => x"fff4b408",
   716 => x"51a08091",
   717 => x"be2d83ff",
   718 => x"e0800883",
   719 => x"fff4b40c",
   720 => x"84801581",
   721 => x"17575576",
   722 => x"7624ffa4",
   723 => x"38a08096",
   724 => x"dd0483ff",
   725 => x"e0800854",
   726 => x"a08096df",
   727 => x"04815473",
   728 => x"83ffe080",
   729 => x"0c029c05",
   730 => x"0d0483ff",
   731 => x"e08c0802",
   732 => x"83ffe08c",
   733 => x"0cff3d0d",
   734 => x"800b83ff",
   735 => x"e08c08fc",
   736 => x"050c83ff",
   737 => x"e08c0888",
   738 => x"05088106",
   739 => x"ff117009",
   740 => x"7083ffe0",
   741 => x"8c088c05",
   742 => x"080683ff",
   743 => x"e08c08fc",
   744 => x"05081183",
   745 => x"ffe08c08",
   746 => x"fc050c83",
   747 => x"ffe08c08",
   748 => x"88050881",
   749 => x"2a83ffe0",
   750 => x"8c088805",
   751 => x"0c83ffe0",
   752 => x"8c088c05",
   753 => x"081083ff",
   754 => x"e08c088c",
   755 => x"050c5151",
   756 => x"515183ff",
   757 => x"e08c0888",
   758 => x"0508802e",
   759 => x"8438ffa2",
   760 => x"3983ffe0",
   761 => x"8c08fc05",
   762 => x"087083ff",
   763 => x"e0800c51",
   764 => x"833d0d83",
   765 => x"ffe08c0c",
   766 => x"04000000",
   767 => x"00ffffff",
   768 => x"ff00ffff",
   769 => x"ffff00ff",
   770 => x"ffffff00",
   771 => x"4d414e49",
   772 => x"46455354",
   773 => x"4d535400",
   774 => x"46415431",
   775 => x"36202020",
   776 => x"00000000",
   777 => x"46415433",
   778 => x"32202020",
   779 => x"00000000",
	others => x"00000000"
);

begin

process (clk)
begin
	if (clk'event and clk = '1') then
		if (from_zpu.memAWriteEnable = '1') and (from_zpu.memBWriteEnable = '1') and (from_zpu.memAAddr=from_zpu.memBAddr) and (from_zpu.memAWrite/=from_zpu.memBWrite) then
			report "write collision" severity failure;
		end if;
	
		if (from_zpu.memAWriteEnable = '1') then
			ram(to_integer(unsigned(from_zpu.memAAddr(maxAddrBit downto 2)))) := from_zpu.memAWrite;
			to_zpu.memARead <= from_zpu.memAWrite;
		else
			to_zpu.memARead <= ram(to_integer(unsigned(from_zpu.memAAddr(maxAddrBit downto 2))));
		end if;
	end if;
end process;

process (clk)
begin
	if (clk'event and clk = '1') then
		if (from_zpu.memBWriteEnable = '1') then
			ram(to_integer(unsigned(from_zpu.memBAddr(maxAddrBit downto 2)))) := from_zpu.memBWrite;
			to_zpu.memBRead <= from_zpu.memBWrite;
		else
			to_zpu.memBRead <= ram(to_integer(unsigned(from_zpu.memBAddr(maxAddrBit downto 2))));
		end if;
	end if;
end process;


end arch;

