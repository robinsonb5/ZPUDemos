-- ZPU
--
-- Copyright 2004-2008 oharboe - �yvind Harboe - oyvind.harboe@zylin.com
-- Modified by Alastair M. Robinson for the ZPUFlex project.
--
-- The FreeBSD license
-- 
-- Redistribution and use in source and binary forms, with or without
-- modification, are permitted provided that the following conditions
-- are met:
-- 
-- 1. Redistributions of source code must retain the above copyright
--    notice, this list of conditions and the following disclaimer.
-- 2. Redistributions in binary form must reproduce the above
--    copyright notice, this list of conditions and the following
--    disclaimer in the documentation and/or other materials
--    provided with the distribution.
-- 
-- THIS SOFTWARE IS PROVIDED BY THE ZPU PROJECT ``AS IS'' AND ANY
-- EXPRESS OR IMPLIED WARRANTIES, INCLUDING, BUT NOT LIMITED TO,
-- THE IMPLIED WARRANTIES OF MERCHANTABILITY AND FITNESS FOR A
-- PARTICULAR PURPOSE ARE DISCLAIMED. IN NO EVENT SHALL THE
-- ZPU PROJECT OR CONTRIBUTORS BE LIABLE FOR ANY DIRECT,
-- INDIRECT, INCIDENTAL, SPECIAL, EXEMPLARY, OR CONSEQUENTIAL DAMAGES
-- (INCLUDING, BUT NOT LIMITED TO, PROCUREMENT OF SUBSTITUTE GOODS
-- OR SERVICES; LOSS OF USE, DATA, OR PROFITS; OR BUSINESS INTERRUPTION)
-- HOWEVER CAUSED AND ON ANY THEORY OF LIABILITY, WHETHER IN CONTRACT,
-- STRICT LIABILITY, OR TORT (INCLUDING NEGLIGENCE OR OTHERWISE)
-- ARISING IN ANY WAY OUT OF THE USE OF THIS SOFTWARE, EVEN IF
-- ADVISED OF THE POSSIBILITY OF SUCH DAMAGE.
-- 
-- The views and conclusions contained in the software and documentation
-- are those of the authors and should not be interpreted as representing
-- official policies, either expressed or implied, of the ZPU Project.

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;


library work;
use work.zpupkg.all;

entity VGATest_ROM is
generic
	(
		maxAddrBitBRAM : integer := maxAddrBitBRAMLimit -- Specify your actual ROM size to save LEs and unnecessary block RAM usage.
	);
port (
	clk : in std_logic;
	areset : in std_logic := '0';
	from_zpu : in ZPU_ToROM;
	to_zpu : out ZPU_FromROM
);
end VGATest_ROM;

architecture arch of VGATest_ROM is

type ram_type is array(natural range 0 to ((2**(maxAddrBitBRAM+1))/4)-1) of std_logic_vector(wordSize-1 downto 0);

shared variable ram : ram_type :=
(
     0 => x"84808080",
     1 => x"8c0b8480",
     2 => x"8081e004",
     3 => x"00848080",
     4 => x"808c04ff",
     5 => x"0d800404",
     6 => x"40000017",
     7 => x"00000000",
     8 => x"84808099",
     9 => x"a0088480",
    10 => x"8099a408",
    11 => x"84808099",
    12 => x"a8088480",
    13 => x"80809808",
    14 => x"2d848080",
    15 => x"99a80c84",
    16 => x"808099a4",
    17 => x"0c848080",
    18 => x"99a00c04",
    19 => x"00000000",
    20 => x"00000000",
    21 => x"00000000",
    22 => x"00000000",
    23 => x"00000000",
    24 => x"71fd0608",
    25 => x"72830609",
    26 => x"81058205",
    27 => x"832b2a83",
    28 => x"ffff0652",
    29 => x"0471fc06",
    30 => x"08728306",
    31 => x"09810583",
    32 => x"05101010",
    33 => x"2a81ff06",
    34 => x"520471fd",
    35 => x"060883ff",
    36 => x"ff738306",
    37 => x"09810582",
    38 => x"05832b2b",
    39 => x"09067383",
    40 => x"ffff0673",
    41 => x"83060981",
    42 => x"05820583",
    43 => x"2b0b2b07",
    44 => x"72fc060c",
    45 => x"51510471",
    46 => x"fc060884",
    47 => x"80809394",
    48 => x"73830610",
    49 => x"10050806",
    50 => x"7381ff06",
    51 => x"73830609",
    52 => x"81058305",
    53 => x"1010102b",
    54 => x"0772fc06",
    55 => x"0c515104",
    56 => x"84808099",
    57 => x"a0708480",
    58 => x"809ac027",
    59 => x"8e388071",
    60 => x"70840553",
    61 => x"0c848080",
    62 => x"81e50484",
    63 => x"8080808c",
    64 => x"51848080",
    65 => x"86cb0402",
    66 => x"c0050d02",
    67 => x"80c4055b",
    68 => x"80707c70",
    69 => x"84055e08",
    70 => x"725f5f5f",
    71 => x"5a7c7084",
    72 => x"055e0857",
    73 => x"80597698",
    74 => x"2a77882b",
    75 => x"58557480",
    76 => x"2e82e738",
    77 => x"7b802e80",
    78 => x"d338805c",
    79 => x"7480e42e",
    80 => x"81d83874",
    81 => x"80f82e81",
    82 => x"d1387480",
    83 => x"e42e81dc",
    84 => x"387480e4",
    85 => x"2680f138",
    86 => x"7480e32e",
    87 => x"80c838a5",
    88 => x"51848080",
    89 => x"85db2d74",
    90 => x"51848080",
    91 => x"85db2d82",
    92 => x"1a811a5a",
    93 => x"5a837925",
    94 => x"ffac3874",
    95 => x"ff9f387e",
    96 => x"84808099",
    97 => x"a00c0280",
    98 => x"c0050d04",
    99 => x"74a52e09",
   100 => x"81069b38",
   101 => x"810b811a",
   102 => x"5a5c8379",
   103 => x"25ff8738",
   104 => x"84808082",
   105 => x"fb047a84",
   106 => x"1c710857",
   107 => x"5c547451",
   108 => x"84808085",
   109 => x"db2d811a",
   110 => x"811a5a5a",
   111 => x"837925fe",
   112 => x"e5388480",
   113 => x"8082fb04",
   114 => x"7480f32e",
   115 => x"81d93874",
   116 => x"80f82e09",
   117 => x"8106ff87",
   118 => x"387d5380",
   119 => x"587d782e",
   120 => x"81e23887",
   121 => x"56729c2a",
   122 => x"73842b54",
   123 => x"5271802e",
   124 => x"83388158",
   125 => x"b7125471",
   126 => x"89248438",
   127 => x"b0125477",
   128 => x"80ea38ff",
   129 => x"16567580",
   130 => x"25db3881",
   131 => x"19598379",
   132 => x"25fe9338",
   133 => x"84808082",
   134 => x"fb047a84",
   135 => x"1c710840",
   136 => x"5c527480",
   137 => x"e42e0981",
   138 => x"06fea638",
   139 => x"7d538058",
   140 => x"7d782e81",
   141 => x"8f388756",
   142 => x"729c2a73",
   143 => x"842b5452",
   144 => x"71802e83",
   145 => x"388158b7",
   146 => x"12547189",
   147 => x"248438b0",
   148 => x"125477af",
   149 => x"38ff1656",
   150 => x"758025dc",
   151 => x"38811959",
   152 => x"837925fd",
   153 => x"c1388480",
   154 => x"8082fb04",
   155 => x"73518480",
   156 => x"8085db2d",
   157 => x"ff165675",
   158 => x"8025fee9",
   159 => x"38848080",
   160 => x"848b0473",
   161 => x"51848080",
   162 => x"85db2dff",
   163 => x"16567580",
   164 => x"25ffa538",
   165 => x"84808084",
   166 => x"dd047984",
   167 => x"808099a0",
   168 => x"0c0280c0",
   169 => x"050d047a",
   170 => x"841c7108",
   171 => x"535c5384",
   172 => x"80808680",
   173 => x"2d811959",
   174 => x"837925fc",
   175 => x"e9388480",
   176 => x"8082fb04",
   177 => x"b0518480",
   178 => x"8085db2d",
   179 => x"81195983",
   180 => x"7925fcd2",
   181 => x"38848080",
   182 => x"82fb0402",
   183 => x"f8050d73",
   184 => x"52c00870",
   185 => x"882a7081",
   186 => x"06515151",
   187 => x"70802ef1",
   188 => x"3871c00c",
   189 => x"71848080",
   190 => x"99a00c02",
   191 => x"88050d04",
   192 => x"02e8050d",
   193 => x"80785755",
   194 => x"75708405",
   195 => x"57085380",
   196 => x"5472982a",
   197 => x"73882b54",
   198 => x"5271802e",
   199 => x"a238c008",
   200 => x"70882a70",
   201 => x"81065151",
   202 => x"5170802e",
   203 => x"f13871c0",
   204 => x"0c811581",
   205 => x"15555583",
   206 => x"7425d638",
   207 => x"71ca3874",
   208 => x"84808099",
   209 => x"a00c0298",
   210 => x"050d0402",
   211 => x"dc050d80",
   212 => x"52848080",
   213 => x"0bfc800c",
   214 => x"81127055",
   215 => x"59848080",
   216 => x"56805584",
   217 => x"fe538114",
   218 => x"83ffff06",
   219 => x"70777084",
   220 => x"05590cfe",
   221 => x"14545472",
   222 => x"8025eb38",
   223 => x"81155583",
   224 => x"df7525df",
   225 => x"38805780",
   226 => x"5584fe53",
   227 => x"fc8008fe",
   228 => x"14545272",
   229 => x"8025f538",
   230 => x"81155583",
   231 => x"df7525e9",
   232 => x"38811757",
   233 => x"b17725df",
   234 => x"38805875",
   235 => x"55805784",
   236 => x"fe538114",
   237 => x"83ffff06",
   238 => x"70767084",
   239 => x"05580cfe",
   240 => x"14545472",
   241 => x"8025eb38",
   242 => x"81175783",
   243 => x"df7725df",
   244 => x"38811858",
   245 => x"937825d3",
   246 => x"38811952",
   247 => x"80518480",
   248 => x"808fd42d",
   249 => x"84808086",
   250 => x"d80402f4",
   251 => x"050d7476",
   252 => x"52538071",
   253 => x"25903870",
   254 => x"52727084",
   255 => x"055408ff",
   256 => x"13535171",
   257 => x"f438028c",
   258 => x"050d0402",
   259 => x"d4050d7c",
   260 => x"7e5c5881",
   261 => x"0b848080",
   262 => x"93a4585a",
   263 => x"83597608",
   264 => x"780c7708",
   265 => x"77085654",
   266 => x"73752e94",
   267 => x"38770853",
   268 => x"74528480",
   269 => x"8093b451",
   270 => x"84808082",
   271 => x"872d805a",
   272 => x"7756807b",
   273 => x"2590387a",
   274 => x"55757084",
   275 => x"055708ff",
   276 => x"16565474",
   277 => x"f4387708",
   278 => x"77085656",
   279 => x"75752e94",
   280 => x"38770853",
   281 => x"74528480",
   282 => x"8093f451",
   283 => x"84808082",
   284 => x"872d805a",
   285 => x"ff198418",
   286 => x"58597880",
   287 => x"25ff9f38",
   288 => x"79848080",
   289 => x"99a00c02",
   290 => x"ac050d04",
   291 => x"02e4050d",
   292 => x"787a5556",
   293 => x"815785aa",
   294 => x"d5aad576",
   295 => x"0cfad5aa",
   296 => x"d5aa0b8c",
   297 => x"170ccc76",
   298 => x"84808081",
   299 => x"b72db30b",
   300 => x"8f178480",
   301 => x"8081b72d",
   302 => x"75085372",
   303 => x"fce2d5aa",
   304 => x"d52e9238",
   305 => x"75085284",
   306 => x"808094b4",
   307 => x"51848080",
   308 => x"82872d80",
   309 => x"578c1608",
   310 => x"5574fad5",
   311 => x"aad4b32e",
   312 => x"93388c16",
   313 => x"08528480",
   314 => x"8094f051",
   315 => x"84808082",
   316 => x"872d8057",
   317 => x"75558074",
   318 => x"258e3874",
   319 => x"70840556",
   320 => x"08ff1555",
   321 => x"5373f438",
   322 => x"75085473",
   323 => x"fce2d5aa",
   324 => x"d52e9238",
   325 => x"75085284",
   326 => x"808095ac",
   327 => x"51848080",
   328 => x"82872d80",
   329 => x"578c1608",
   330 => x"5372fad5",
   331 => x"aad4b32e",
   332 => x"93388c16",
   333 => x"08528480",
   334 => x"8095e851",
   335 => x"84808082",
   336 => x"872d8057",
   337 => x"76848080",
   338 => x"99a00c02",
   339 => x"9c050d04",
   340 => x"02c4050d",
   341 => x"605b8062",
   342 => x"90808029",
   343 => x"ff058480",
   344 => x"8096a453",
   345 => x"405a8480",
   346 => x"8082872d",
   347 => x"80e1b357",
   348 => x"80fe5eae",
   349 => x"51848080",
   350 => x"85db2d76",
   351 => x"1070962a",
   352 => x"81065657",
   353 => x"74802e85",
   354 => x"38768107",
   355 => x"5776952a",
   356 => x"81065877",
   357 => x"802e8538",
   358 => x"76813257",
   359 => x"7877077f",
   360 => x"06775e59",
   361 => x"8fffff58",
   362 => x"76bfffff",
   363 => x"06707a32",
   364 => x"822b7c11",
   365 => x"5157760c",
   366 => x"76107096",
   367 => x"2a810656",
   368 => x"5774802e",
   369 => x"85387681",
   370 => x"07577695",
   371 => x"2a810655",
   372 => x"74802e85",
   373 => x"38768132",
   374 => x"57ff1858",
   375 => x"778025c8",
   376 => x"387c578f",
   377 => x"ffff5876",
   378 => x"bfffff06",
   379 => x"707a3282",
   380 => x"2b7c0570",
   381 => x"08575e56",
   382 => x"74762e80",
   383 => x"ea38807a",
   384 => x"53848080",
   385 => x"96b4525c",
   386 => x"84808082",
   387 => x"872d7454",
   388 => x"75537552",
   389 => x"84808096",
   390 => x"c8518480",
   391 => x"8082872d",
   392 => x"7b5a7610",
   393 => x"70962a81",
   394 => x"06575775",
   395 => x"802e8538",
   396 => x"76810757",
   397 => x"76952a81",
   398 => x"06557480",
   399 => x"2e853876",
   400 => x"813257ff",
   401 => x"18587780",
   402 => x"25ff9c38",
   403 => x"ff1e5e7d",
   404 => x"fea1388a",
   405 => x"51848080",
   406 => x"85db2d7b",
   407 => x"84808099",
   408 => x"a00c02bc",
   409 => x"050d0481",
   410 => x"1a5a8480",
   411 => x"808ca204",
   412 => x"02cc050d",
   413 => x"7e605e58",
   414 => x"815a805b",
   415 => x"80c07a58",
   416 => x"5c85ada9",
   417 => x"89bb780c",
   418 => x"79598156",
   419 => x"97557676",
   420 => x"07822b78",
   421 => x"11515485",
   422 => x"ada989bb",
   423 => x"740c7510",
   424 => x"ff165656",
   425 => x"748025e6",
   426 => x"38761081",
   427 => x"1a5a5798",
   428 => x"7925d738",
   429 => x"7756807d",
   430 => x"2590387c",
   431 => x"55757084",
   432 => x"055708ff",
   433 => x"16565474",
   434 => x"f4388157",
   435 => x"ff8787a5",
   436 => x"c3780c97",
   437 => x"5976822b",
   438 => x"78117008",
   439 => x"5f56567c",
   440 => x"ff8787a5",
   441 => x"c32e80cc",
   442 => x"38740854",
   443 => x"7385ada9",
   444 => x"89bb2e94",
   445 => x"38807508",
   446 => x"54765384",
   447 => x"808096f0",
   448 => x"525a8480",
   449 => x"8082872d",
   450 => x"7610ff1a",
   451 => x"5a577880",
   452 => x"25c3387a",
   453 => x"822b5675",
   454 => x"b1387b52",
   455 => x"84808097",
   456 => x"90518480",
   457 => x"8082872d",
   458 => x"7b848080",
   459 => x"99a00c02",
   460 => x"b4050d04",
   461 => x"7a770777",
   462 => x"10ff1b5b",
   463 => x"585b7880",
   464 => x"25ff9238",
   465 => x"8480808e",
   466 => x"93047552",
   467 => x"84808097",
   468 => x"cc518480",
   469 => x"8082872d",
   470 => x"75992a81",
   471 => x"32810670",
   472 => x"09810571",
   473 => x"07700970",
   474 => x"9f2c7d06",
   475 => x"79109fff",
   476 => x"fffc0660",
   477 => x"812a415a",
   478 => x"5d575859",
   479 => x"75da3879",
   480 => x"09810570",
   481 => x"7b079f2a",
   482 => x"55567bbf",
   483 => x"26843873",
   484 => x"9d388170",
   485 => x"53848080",
   486 => x"9790525c",
   487 => x"84808082",
   488 => x"872d7b84",
   489 => x"808099a0",
   490 => x"0c02b405",
   491 => x"0d048480",
   492 => x"8097e451",
   493 => x"84808082",
   494 => x"872d7b52",
   495 => x"84808097",
   496 => x"90518480",
   497 => x"8082872d",
   498 => x"7b848080",
   499 => x"99a00c02",
   500 => x"b4050d04",
   501 => x"02d4050d",
   502 => x"7c578170",
   503 => x"84808093",
   504 => x"a45b595b",
   505 => x"835a7808",
   506 => x"770c7608",
   507 => x"79085654",
   508 => x"73752e94",
   509 => x"38760853",
   510 => x"74528480",
   511 => x"8093b451",
   512 => x"84808082",
   513 => x"872d8058",
   514 => x"76569fff",
   515 => x"55757084",
   516 => x"055708ff",
   517 => x"16565474",
   518 => x"8025f238",
   519 => x"76087908",
   520 => x"56567575",
   521 => x"2e943876",
   522 => x"08537452",
   523 => x"84808093",
   524 => x"f4518480",
   525 => x"8082872d",
   526 => x"8058ff1a",
   527 => x"841a5a5a",
   528 => x"798025ff",
   529 => x"a1387781",
   530 => x"fd38775b",
   531 => x"815885aa",
   532 => x"d5aad577",
   533 => x"0cfad5aa",
   534 => x"d5aa0b8c",
   535 => x"180ccc77",
   536 => x"84808081",
   537 => x"b72db30b",
   538 => x"8f188480",
   539 => x"8081b72d",
   540 => x"76085574",
   541 => x"fce2d5aa",
   542 => x"d52e9238",
   543 => x"76085284",
   544 => x"808094b4",
   545 => x"51848080",
   546 => x"82872d80",
   547 => x"588c1708",
   548 => x"5978fad5",
   549 => x"aad4b32e",
   550 => x"93388c17",
   551 => x"08528480",
   552 => x"8094f051",
   553 => x"84808082",
   554 => x"872d8058",
   555 => x"76569fff",
   556 => x"55757084",
   557 => x"055708ff",
   558 => x"16565474",
   559 => x"8025f238",
   560 => x"76085a79",
   561 => x"fce2d5aa",
   562 => x"d52e9238",
   563 => x"76085284",
   564 => x"808095ac",
   565 => x"51848080",
   566 => x"82872d80",
   567 => x"588c1708",
   568 => x"5473fad5",
   569 => x"aad4b32e",
   570 => x"80ee388c",
   571 => x"17085284",
   572 => x"808095e8",
   573 => x"51848080",
   574 => x"82872d80",
   575 => x"58775ba0",
   576 => x"80527651",
   577 => x"8480808c",
   578 => x"f02d8480",
   579 => x"8099a008",
   580 => x"54848080",
   581 => x"99a00880",
   582 => x"e9388480",
   583 => x"8099a008",
   584 => x"5b735276",
   585 => x"51848080",
   586 => x"8ad02d84",
   587 => x"808099a0",
   588 => x"08be3884",
   589 => x"808099a0",
   590 => x"085b7a84",
   591 => x"808099a0",
   592 => x"0c02ac05",
   593 => x"0d048480",
   594 => x"8098b051",
   595 => x"84808082",
   596 => x"872d8480",
   597 => x"8090cc04",
   598 => x"77802eff",
   599 => x"a0388480",
   600 => x"8098d451",
   601 => x"84808082",
   602 => x"872d8480",
   603 => x"8091ff04",
   604 => x"84808098",
   605 => x"f0518480",
   606 => x"8082872d",
   607 => x"84808092",
   608 => x"ba048480",
   609 => x"80998851",
   610 => x"84808082",
   611 => x"872d8480",
   612 => x"8092a104",
   613 => x"00ffffff",
   614 => x"ff00ffff",
   615 => x"ffff00ff",
   616 => x"ffffff00",
   617 => x"00000000",
   618 => x"55555555",
   619 => x"aaaaaaaa",
   620 => x"ffffffff",
   621 => x"53616e69",
   622 => x"74792063",
   623 => x"6865636b",
   624 => x"20666169",
   625 => x"6c656420",
   626 => x"28626566",
   627 => x"6f726520",
   628 => x"63616368",
   629 => x"65207265",
   630 => x"66726573",
   631 => x"6829206f",
   632 => x"6e203078",
   633 => x"25642028",
   634 => x"676f7420",
   635 => x"30782564",
   636 => x"290a0000",
   637 => x"53616e69",
   638 => x"74792063",
   639 => x"6865636b",
   640 => x"20666169",
   641 => x"6c656420",
   642 => x"28616674",
   643 => x"65722063",
   644 => x"61636865",
   645 => x"20726566",
   646 => x"72657368",
   647 => x"29206f6e",
   648 => x"20307825",
   649 => x"64202867",
   650 => x"6f742030",
   651 => x"78256429",
   652 => x"0a000000",
   653 => x"42797465",
   654 => x"20636865",
   655 => x"636b2066",
   656 => x"61696c65",
   657 => x"64202862",
   658 => x"65666f72",
   659 => x"65206361",
   660 => x"63686520",
   661 => x"72656672",
   662 => x"65736829",
   663 => x"20617420",
   664 => x"30202867",
   665 => x"6f742030",
   666 => x"78256429",
   667 => x"0a000000",
   668 => x"42797465",
   669 => x"20636865",
   670 => x"636b2066",
   671 => x"61696c65",
   672 => x"64202862",
   673 => x"65666f72",
   674 => x"65206361",
   675 => x"63686520",
   676 => x"72656672",
   677 => x"65736829",
   678 => x"20617420",
   679 => x"33202867",
   680 => x"6f742030",
   681 => x"78256429",
   682 => x"0a000000",
   683 => x"42797465",
   684 => x"20636865",
   685 => x"636b2066",
   686 => x"61696c65",
   687 => x"64202861",
   688 => x"66746572",
   689 => x"20636163",
   690 => x"68652072",
   691 => x"65667265",
   692 => x"73682920",
   693 => x"61742030",
   694 => x"2028676f",
   695 => x"74203078",
   696 => x"2564290a",
   697 => x"00000000",
   698 => x"42797465",
   699 => x"20636865",
   700 => x"636b2066",
   701 => x"61696c65",
   702 => x"64202861",
   703 => x"66746572",
   704 => x"20636163",
   705 => x"68652072",
   706 => x"65667265",
   707 => x"73682920",
   708 => x"61742033",
   709 => x"2028676f",
   710 => x"74203078",
   711 => x"2564290a",
   712 => x"00000000",
   713 => x"43686563",
   714 => x"6b696e67",
   715 => x"206d656d",
   716 => x"6f727900",
   717 => x"30782564",
   718 => x"20676f6f",
   719 => x"64207265",
   720 => x"6164732c",
   721 => x"20000000",
   722 => x"4572726f",
   723 => x"72206174",
   724 => x"20307825",
   725 => x"642c2065",
   726 => x"78706563",
   727 => x"74656420",
   728 => x"30782564",
   729 => x"2c20676f",
   730 => x"74203078",
   731 => x"25640a00",
   732 => x"42616420",
   733 => x"64617461",
   734 => x"20666f75",
   735 => x"6e642061",
   736 => x"74203078",
   737 => x"25642028",
   738 => x"30782564",
   739 => x"290a0000",
   740 => x"53445241",
   741 => x"4d207369",
   742 => x"7a652028",
   743 => x"61737375",
   744 => x"6d696e67",
   745 => x"206e6f20",
   746 => x"61646472",
   747 => x"65737320",
   748 => x"6661756c",
   749 => x"74732920",
   750 => x"69732030",
   751 => x"78256420",
   752 => x"6d656761",
   753 => x"62797465",
   754 => x"730a0000",
   755 => x"416c6961",
   756 => x"73657320",
   757 => x"666f756e",
   758 => x"64206174",
   759 => x"20307825",
   760 => x"640a0000",
   761 => x"28416c69",
   762 => x"61736573",
   763 => x"2070726f",
   764 => x"6261626c",
   765 => x"79207369",
   766 => x"6d706c79",
   767 => x"20696e64",
   768 => x"69636174",
   769 => x"65207468",
   770 => x"61742052",
   771 => x"414d0a69",
   772 => x"7320736d",
   773 => x"616c6c65",
   774 => x"72207468",
   775 => x"616e2036",
   776 => x"34206d65",
   777 => x"67616279",
   778 => x"74657329",
   779 => x"0a000000",
   780 => x"46697273",
   781 => x"74207374",
   782 => x"61676520",
   783 => x"73616e69",
   784 => x"74792063",
   785 => x"6865636b",
   786 => x"20706173",
   787 => x"7365642e",
   788 => x"0a000000",
   789 => x"42797465",
   790 => x"20286471",
   791 => x"6d292063",
   792 => x"6865636b",
   793 => x"20706173",
   794 => x"7365640a",
   795 => x"00000000",
   796 => x"4c465352",
   797 => x"20636865",
   798 => x"636b2070",
   799 => x"61737365",
   800 => x"642e0a0a",
   801 => x"00000000",
   802 => x"41646472",
   803 => x"65737320",
   804 => x"63686563",
   805 => x"6b207061",
   806 => x"73736564",
   807 => x"2e0a0000",
	others => x"00000000"
);

begin

process (clk)
begin
	if (clk'event and clk = '1') then
		if (from_zpu.memAWriteEnable = '1') and (from_zpu.memBWriteEnable = '1') and (from_zpu.memAAddr=from_zpu.memBAddr) and (from_zpu.memAWrite/=from_zpu.memBWrite) then
			report "write collision" severity failure;
		end if;
	
		if (from_zpu.memAWriteEnable = '1') then
			ram(to_integer(unsigned(from_zpu.memAAddr(maxAddrBitBRAM downto 2)))) := from_zpu.memAWrite;
			to_zpu.memARead <= from_zpu.memAWrite;
		else
			to_zpu.memARead <= ram(to_integer(unsigned(from_zpu.memAAddr(maxAddrBitBRAM downto 2))));
		end if;
	end if;
end process;

process (clk)
begin
	if (clk'event and clk = '1') then
		if (from_zpu.memBWriteEnable = '1') then
			ram(to_integer(unsigned(from_zpu.memBAddr(maxAddrBitBRAM downto 2)))) := from_zpu.memBWrite;
			to_zpu.memBRead <= from_zpu.memBWrite;
		else
			to_zpu.memBRead <= ram(to_integer(unsigned(from_zpu.memBAddr(maxAddrBitBRAM downto 2))));
		end if;
	end if;
end process;


end arch;

