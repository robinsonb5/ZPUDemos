-- ZPU
--
-- Copyright 2004-2008 oharboe - �yvind Harboe - oyvind.harboe@zylin.com
-- Modified by Alastair M. Robinson for the ZPUFlex project.
--
-- The FreeBSD license
-- 
-- Redistribution and use in source and binary forms, with or without
-- modification, are permitted provided that the following conditions
-- are met:
-- 
-- 1. Redistributions of source code must retain the above copyright
--    notice, this list of conditions and the following disclaimer.
-- 2. Redistributions in binary form must reproduce the above
--    copyright notice, this list of conditions and the following
--    disclaimer in the documentation and/or other materials
--    provided with the distribution.
-- 
-- THIS SOFTWARE IS PROVIDED BY THE ZPU PROJECT ``AS IS'' AND ANY
-- EXPRESS OR IMPLIED WARRANTIES, INCLUDING, BUT NOT LIMITED TO,
-- THE IMPLIED WARRANTIES OF MERCHANTABILITY AND FITNESS FOR A
-- PARTICULAR PURPOSE ARE DISCLAIMED. IN NO EVENT SHALL THE
-- ZPU PROJECT OR CONTRIBUTORS BE LIABLE FOR ANY DIRECT,
-- INDIRECT, INCIDENTAL, SPECIAL, EXEMPLARY, OR CONSEQUENTIAL DAMAGES
-- (INCLUDING, BUT NOT LIMITED TO, PROCUREMENT OF SUBSTITUTE GOODS
-- OR SERVICES; LOSS OF USE, DATA, OR PROFITS; OR BUSINESS INTERRUPTION)
-- HOWEVER CAUSED AND ON ANY THEORY OF LIABILITY, WHETHER IN CONTRACT,
-- STRICT LIABILITY, OR TORT (INCLUDING NEGLIGENCE OR OTHERWISE)
-- ARISING IN ANY WAY OUT OF THE USE OF THIS SOFTWARE, EVEN IF
-- ADVISED OF THE POSSIBILITY OF SUCH DAMAGE.
-- 
-- The views and conclusions contained in the software and documentation
-- are those of the authors and should not be interpreted as representing
-- official policies, either expressed or implied, of the ZPU Project.

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;


library work;
use work.zpu_config.all;
use work.zpupkg.all;

entity Dhrystone_fast_ROM is
generic
	(
		maxAddrBit : integer := maxAddrBitBRAMLimit -- Specify your actual ROM size to save LEs and unnecessary block RAM usage.
	);
port (
	clk : in std_logic;
	areset : in std_logic := '0';
	from_zpu : in ZPU_ToROM;
	to_zpu : out ZPU_FromROM
);
end Dhrystone_fast_ROM;

architecture arch of Dhrystone_fast_ROM is

type ram_type is array(natural range 0 to ((2**(maxAddrBit+1))/4)-1) of std_logic_vector(wordSize-1 downto 0);

shared variable ram : ram_type :=
(
     0 => x"0b0b0b88",
     1 => x"dd040000",
     2 => x"00000000",
     3 => x"00000000",
     4 => x"00000000",
     5 => x"00000000",
     6 => x"00000000",
     7 => x"00000000",
     8 => x"04000000",
     9 => x"00000000",
    10 => x"00000000",
    11 => x"00000000",
    12 => x"00000000",
    13 => x"00000000",
    14 => x"00000000",
    15 => x"00000000",
    16 => x"71fd0608",
    17 => x"72830609",
    18 => x"81058205",
    19 => x"832b2a83",
    20 => x"ffff0652",
    21 => x"04000000",
    22 => x"00000000",
    23 => x"00000000",
    24 => x"71fd0608",
    25 => x"83ffff73",
    26 => x"83060981",
    27 => x"05820583",
    28 => x"2b2b0906",
    29 => x"7383ffff",
    30 => x"0b0b0b0b",
    31 => x"83a50400",
    32 => x"72098105",
    33 => x"72057373",
    34 => x"09060906",
    35 => x"73097306",
    36 => x"070a8106",
    37 => x"53510400",
    38 => x"00000000",
    39 => x"00000000",
    40 => x"72722473",
    41 => x"732e0753",
    42 => x"51040000",
    43 => x"00000000",
    44 => x"00000000",
    45 => x"00000000",
    46 => x"00000000",
    47 => x"00000000",
    48 => x"71737109",
    49 => x"71068106",
    50 => x"09810572",
    51 => x"0a100a72",
    52 => x"0a100a31",
    53 => x"050a8106",
    54 => x"51515351",
    55 => x"04000000",
    56 => x"72722673",
    57 => x"732e0753",
    58 => x"51040000",
    59 => x"00000000",
    60 => x"00000000",
    61 => x"00000000",
    62 => x"00000000",
    63 => x"00000000",
    64 => x"00000000",
    65 => x"00000000",
    66 => x"00000000",
    67 => x"00000000",
    68 => x"00000000",
    69 => x"00000000",
    70 => x"00000000",
    71 => x"00000000",
    72 => x"0b0b0b88",
    73 => x"ba040000",
    74 => x"00000000",
    75 => x"00000000",
    76 => x"00000000",
    77 => x"00000000",
    78 => x"00000000",
    79 => x"00000000",
    80 => x"720a722b",
    81 => x"0a535104",
    82 => x"00000000",
    83 => x"00000000",
    84 => x"00000000",
    85 => x"00000000",
    86 => x"00000000",
    87 => x"00000000",
    88 => x"72729f06",
    89 => x"0981050b",
    90 => x"0b0b889f",
    91 => x"05040000",
    92 => x"00000000",
    93 => x"00000000",
    94 => x"00000000",
    95 => x"00000000",
    96 => x"72722aff",
    97 => x"739f062a",
    98 => x"0974090a",
    99 => x"8106ff05",
   100 => x"06075351",
   101 => x"04000000",
   102 => x"00000000",
   103 => x"00000000",
   104 => x"71715351",
   105 => x"04067383",
   106 => x"06098105",
   107 => x"8205832b",
   108 => x"0b2b0772",
   109 => x"fc060c51",
   110 => x"51040000",
   111 => x"00000000",
   112 => x"72098105",
   113 => x"72050970",
   114 => x"81050906",
   115 => x"0a810653",
   116 => x"51040000",
   117 => x"00000000",
   118 => x"00000000",
   119 => x"00000000",
   120 => x"72098105",
   121 => x"72050970",
   122 => x"81050906",
   123 => x"0a098106",
   124 => x"53510400",
   125 => x"00000000",
   126 => x"00000000",
   127 => x"00000000",
   128 => x"71098105",
   129 => x"52040000",
   130 => x"00000000",
   131 => x"00000000",
   132 => x"00000000",
   133 => x"00000000",
   134 => x"00000000",
   135 => x"00000000",
   136 => x"72720981",
   137 => x"05055351",
   138 => x"04000000",
   139 => x"00000000",
   140 => x"00000000",
   141 => x"00000000",
   142 => x"00000000",
   143 => x"00000000",
   144 => x"72097206",
   145 => x"73730906",
   146 => x"07535104",
   147 => x"00000000",
   148 => x"00000000",
   149 => x"00000000",
   150 => x"00000000",
   151 => x"00000000",
   152 => x"71fc0608",
   153 => x"72830609",
   154 => x"81058305",
   155 => x"1010102a",
   156 => x"81ff0652",
   157 => x"04000000",
   158 => x"00000000",
   159 => x"00000000",
   160 => x"71fc0608",
   161 => x"0b0b0ba1",
   162 => x"8c738306",
   163 => x"10100508",
   164 => x"060b0b0b",
   165 => x"88a20400",
   166 => x"00000000",
   167 => x"00000000",
   168 => x"88088c08",
   169 => x"90087575",
   170 => x"0b0b0b99",
   171 => x"ff2d5050",
   172 => x"88085690",
   173 => x"0c8c0c88",
   174 => x"0c510400",
   175 => x"00000000",
   176 => x"88088c08",
   177 => x"90087575",
   178 => x"0b0b0b9b",
   179 => x"b12d5050",
   180 => x"88085690",
   181 => x"0c8c0c88",
   182 => x"0c510400",
   183 => x"00000000",
   184 => x"72097081",
   185 => x"0509060a",
   186 => x"8106ff05",
   187 => x"70547106",
   188 => x"73097274",
   189 => x"05ff0506",
   190 => x"07515151",
   191 => x"04000000",
   192 => x"72097081",
   193 => x"0509060a",
   194 => x"098106ff",
   195 => x"05705471",
   196 => x"06730972",
   197 => x"7405ff05",
   198 => x"06075151",
   199 => x"51040000",
   200 => x"05ff0504",
   201 => x"00000000",
   202 => x"00000000",
   203 => x"00000000",
   204 => x"00000000",
   205 => x"00000000",
   206 => x"00000000",
   207 => x"00000000",
   208 => x"04000000",
   209 => x"00000000",
   210 => x"00000000",
   211 => x"00000000",
   212 => x"00000000",
   213 => x"00000000",
   214 => x"00000000",
   215 => x"00000000",
   216 => x"71810552",
   217 => x"04000000",
   218 => x"00000000",
   219 => x"00000000",
   220 => x"00000000",
   221 => x"00000000",
   222 => x"00000000",
   223 => x"00000000",
   224 => x"00000000",
   225 => x"00000000",
   226 => x"00000000",
   227 => x"00000000",
   228 => x"00000000",
   229 => x"00000000",
   230 => x"00000000",
   231 => x"00000000",
   232 => x"02840572",
   233 => x"10100552",
   234 => x"04000000",
   235 => x"00000000",
   236 => x"00000000",
   237 => x"00000000",
   238 => x"00000000",
   239 => x"00000000",
   240 => x"00000000",
   241 => x"00000000",
   242 => x"00000000",
   243 => x"00000000",
   244 => x"00000000",
   245 => x"00000000",
   246 => x"00000000",
   247 => x"00000000",
   248 => x"717105ff",
   249 => x"05715351",
   250 => x"020d0400",
   251 => x"00000000",
   252 => x"00000000",
   253 => x"00000000",
   254 => x"00000000",
   255 => x"00000000",
   256 => x"10101010",
   257 => x"10101010",
   258 => x"10101010",
   259 => x"10101010",
   260 => x"10101010",
   261 => x"10101010",
   262 => x"10101010",
   263 => x"10101053",
   264 => x"51047381",
   265 => x"ff067383",
   266 => x"06098105",
   267 => x"83051010",
   268 => x"102b0772",
   269 => x"fc060c51",
   270 => x"51047272",
   271 => x"80728106",
   272 => x"ff050972",
   273 => x"06057110",
   274 => x"52720a10",
   275 => x"0a5372ed",
   276 => x"38515153",
   277 => x"51040000",
   278 => x"800488da",
   279 => x"0488da0b",
   280 => x"8fad0402",
   281 => x"c0050d02",
   282 => x"80c4050b",
   283 => x"0b0ba6b4",
   284 => x"5a5c807c",
   285 => x"7084055e",
   286 => x"08715f5f",
   287 => x"577d7084",
   288 => x"055f0856",
   289 => x"80587598",
   290 => x"2a76882b",
   291 => x"57557480",
   292 => x"2e82d038",
   293 => x"7c802eb9",
   294 => x"38805d74",
   295 => x"80e42e81",
   296 => x"9f387480",
   297 => x"e42680dc",
   298 => x"387480e3",
   299 => x"2eba38a5",
   300 => x"518bec2d",
   301 => x"74518bec",
   302 => x"2d821757",
   303 => x"81185883",
   304 => x"7825c338",
   305 => x"74ffb638",
   306 => x"7e880c02",
   307 => x"80c0050d",
   308 => x"0474a52e",
   309 => x"09810698",
   310 => x"38810b81",
   311 => x"19595d83",
   312 => x"7825ffa2",
   313 => x"3889c404",
   314 => x"7b841d71",
   315 => x"08575d5a",
   316 => x"74518bec",
   317 => x"2d811781",
   318 => x"19595783",
   319 => x"7825ff86",
   320 => x"3889c404",
   321 => x"7480f32e",
   322 => x"098106ff",
   323 => x"a2387b84",
   324 => x"1d710870",
   325 => x"545b5d54",
   326 => x"8c8d2d80",
   327 => x"0bff1155",
   328 => x"53807325",
   329 => x"ff963878",
   330 => x"7081055a",
   331 => x"84e02d70",
   332 => x"52558bec",
   333 => x"2d811774",
   334 => x"ff165654",
   335 => x"578aa104",
   336 => x"7b841d71",
   337 => x"080b0b0b",
   338 => x"a6b40b0b",
   339 => x"0b0ba5e4",
   340 => x"615f585e",
   341 => x"525d5372",
   342 => x"ba38b00b",
   343 => x"0b0b0ba5",
   344 => x"e40b8580",
   345 => x"2d811454",
   346 => x"ff145473",
   347 => x"84e02d7b",
   348 => x"7081055d",
   349 => x"85802d81",
   350 => x"1a5a730b",
   351 => x"0b0ba5e4",
   352 => x"2e098106",
   353 => x"e338807b",
   354 => x"85802d79",
   355 => x"ff115553",
   356 => x"8aa1048a",
   357 => x"52725199",
   358 => x"da2d8808",
   359 => x"0b0b0ba1",
   360 => x"9c0584e0",
   361 => x"2d747081",
   362 => x"05568580",
   363 => x"2d8a5272",
   364 => x"5199b52d",
   365 => x"88085388",
   366 => x"08d93873",
   367 => x"0b0b0ba5",
   368 => x"e42ec338",
   369 => x"ff145473",
   370 => x"84e02d7b",
   371 => x"7081055d",
   372 => x"85802d81",
   373 => x"1a5a730b",
   374 => x"0b0ba5e4",
   375 => x"2effa738",
   376 => x"8ae80476",
   377 => x"880c0280",
   378 => x"c0050d04",
   379 => x"02f8050d",
   380 => x"7352c008",
   381 => x"70882a70",
   382 => x"81065151",
   383 => x"5170802e",
   384 => x"f13871c0",
   385 => x"0c71880c",
   386 => x"0288050d",
   387 => x"0402e805",
   388 => x"0d775675",
   389 => x"70840557",
   390 => x"08538054",
   391 => x"72982a73",
   392 => x"882b5452",
   393 => x"71802ea2",
   394 => x"38c00870",
   395 => x"882a7081",
   396 => x"06515151",
   397 => x"70802ef1",
   398 => x"3871c00c",
   399 => x"81158115",
   400 => x"55558374",
   401 => x"25d63871",
   402 => x"ca387488",
   403 => x"0c029805",
   404 => x"0d04c808",
   405 => x"880c0402",
   406 => x"fc050d80",
   407 => x"c10b80f6",
   408 => x"800b8580",
   409 => x"2d800b80",
   410 => x"f8980c70",
   411 => x"880c0284",
   412 => x"050d0402",
   413 => x"f8050d80",
   414 => x"0b80f680",
   415 => x"0b84e02d",
   416 => x"52527080",
   417 => x"c12e9d38",
   418 => x"7180f898",
   419 => x"080780f8",
   420 => x"980c80c2",
   421 => x"0b80f684",
   422 => x"0b85802d",
   423 => x"70880c02",
   424 => x"88050d04",
   425 => x"810b80f8",
   426 => x"98080780",
   427 => x"f8980c80",
   428 => x"c20b80f6",
   429 => x"840b8580",
   430 => x"2d70880c",
   431 => x"0288050d",
   432 => x"0402f005",
   433 => x"0d757008",
   434 => x"8a055353",
   435 => x"80f6800b",
   436 => x"84e02d51",
   437 => x"7080c12e",
   438 => x"8c3873f0",
   439 => x"3870880c",
   440 => x"0290050d",
   441 => x"04ff1270",
   442 => x"80f5fc08",
   443 => x"31740c88",
   444 => x"0c029005",
   445 => x"0d0402ec",
   446 => x"050d80f6",
   447 => x"a8085574",
   448 => x"802e8c38",
   449 => x"76750871",
   450 => x"0c80f6a8",
   451 => x"0856548c",
   452 => x"155380f5",
   453 => x"fc08528a",
   454 => x"51978b2d",
   455 => x"73880c02",
   456 => x"94050d04",
   457 => x"02e8050d",
   458 => x"77700856",
   459 => x"56b05380",
   460 => x"f6a80852",
   461 => x"74519edd",
   462 => x"2d850b8c",
   463 => x"170c850b",
   464 => x"8c160c75",
   465 => x"08750c80",
   466 => x"f6a80854",
   467 => x"73802e8a",
   468 => x"38730875",
   469 => x"0c80f6a8",
   470 => x"08548c14",
   471 => x"5380f5fc",
   472 => x"08528a51",
   473 => x"978b2d84",
   474 => x"1508ae38",
   475 => x"860b8c16",
   476 => x"0c881552",
   477 => x"88160851",
   478 => x"96a52d80",
   479 => x"f6a80870",
   480 => x"08760c54",
   481 => x"8c157054",
   482 => x"548a5273",
   483 => x"0851978b",
   484 => x"2d73880c",
   485 => x"0298050d",
   486 => x"04750854",
   487 => x"b0537352",
   488 => x"75519edd",
   489 => x"2d73880c",
   490 => x"0298050d",
   491 => x"0402c805",
   492 => x"0d80f594",
   493 => x"0b80f5c8",
   494 => x"0c80f5cc",
   495 => x"0b80f6a8",
   496 => x"0c80f594",
   497 => x"0b80f5cc",
   498 => x"0c800b80",
   499 => x"f5cc0b84",
   500 => x"050c820b",
   501 => x"80f5cc0b",
   502 => x"88050ca8",
   503 => x"0b80f5cc",
   504 => x"0b8c050c",
   505 => x"9f53a1b0",
   506 => x"5280f5dc",
   507 => x"519edd2d",
   508 => x"9f53a1d0",
   509 => x"5280f7f8",
   510 => x"519edd2d",
   511 => x"8a0bb3e0",
   512 => x"0ca4b051",
   513 => x"88e32da1",
   514 => x"f05188e3",
   515 => x"2da4b051",
   516 => x"88e32da5",
   517 => x"e008802e",
   518 => x"849138a2",
   519 => x"a05188e3",
   520 => x"2da4b051",
   521 => x"88e32da5",
   522 => x"dc0852a2",
   523 => x"cc5188e3",
   524 => x"2dc80870",
   525 => x"a7800c56",
   526 => x"8158800b",
   527 => x"a5dc0825",
   528 => x"82dc3802",
   529 => x"ac055b80",
   530 => x"c10b80f6",
   531 => x"800b8580",
   532 => x"2d810b80",
   533 => x"f8980c80",
   534 => x"c20b80f6",
   535 => x"840b8580",
   536 => x"2d825c83",
   537 => x"5a9f53a2",
   538 => x"fc5280f6",
   539 => x"88519edd",
   540 => x"2d815d80",
   541 => x"0b80f688",
   542 => x"5380f7f8",
   543 => x"525598bd",
   544 => x"2d880875",
   545 => x"2e098106",
   546 => x"83388155",
   547 => x"7480f898",
   548 => x"0c7b7057",
   549 => x"55748325",
   550 => x"a1387410",
   551 => x"1015fd05",
   552 => x"5e02b805",
   553 => x"fc055383",
   554 => x"52755197",
   555 => x"8b2d811c",
   556 => x"705d7057",
   557 => x"55837524",
   558 => x"e1387d54",
   559 => x"7453a784",
   560 => x"5280f6b0",
   561 => x"51979d2d",
   562 => x"80f6a808",
   563 => x"70085757",
   564 => x"b0537652",
   565 => x"75519edd",
   566 => x"2d850b8c",
   567 => x"180c850b",
   568 => x"8c170c76",
   569 => x"08760c80",
   570 => x"f6a80855",
   571 => x"74802e8a",
   572 => x"38740876",
   573 => x"0c80f6a8",
   574 => x"08558c15",
   575 => x"5380f5fc",
   576 => x"08528a51",
   577 => x"978b2d84",
   578 => x"160883d8",
   579 => x"38860b8c",
   580 => x"170c8816",
   581 => x"52881708",
   582 => x"5196a52d",
   583 => x"80f6a808",
   584 => x"7008770c",
   585 => x"578c1670",
   586 => x"54558a52",
   587 => x"74085197",
   588 => x"8b2d80c1",
   589 => x"0b80f684",
   590 => x"0b84e02d",
   591 => x"56567575",
   592 => x"26a53880",
   593 => x"c3527551",
   594 => x"98892d88",
   595 => x"087d2e82",
   596 => x"e2388116",
   597 => x"7081ff06",
   598 => x"80f6840b",
   599 => x"84e02d52",
   600 => x"57557476",
   601 => x"27dd3879",
   602 => x"7c297e53",
   603 => x"5199ff2d",
   604 => x"88085c88",
   605 => x"088a0580",
   606 => x"f6800b84",
   607 => x"e02d80f5",
   608 => x"fc085957",
   609 => x"557580c1",
   610 => x"2e82f438",
   611 => x"78f73881",
   612 => x"1858a5dc",
   613 => x"087825fd",
   614 => x"ae38a780",
   615 => x"0856c808",
   616 => x"7080f5c4",
   617 => x"0c707731",
   618 => x"70a6fc0c",
   619 => x"53a39c52",
   620 => x"5b88e32d",
   621 => x"a6fc0856",
   622 => x"80f77625",
   623 => x"80f338a5",
   624 => x"dc087053",
   625 => x"7687e829",
   626 => x"525a99ff",
   627 => x"2d8808a6",
   628 => x"f40c7552",
   629 => x"7987e829",
   630 => x"5199ff2d",
   631 => x"8808a6f8",
   632 => x"0c755279",
   633 => x"84b92951",
   634 => x"99ff2d88",
   635 => x"0880f6ac",
   636 => x"0ca3ac51",
   637 => x"88e32da6",
   638 => x"f40852a3",
   639 => x"dc5188e3",
   640 => x"2da3e451",
   641 => x"88e32da6",
   642 => x"f80852a3",
   643 => x"dc5188e3",
   644 => x"2d80f6ac",
   645 => x"0852a494",
   646 => x"5188e32d",
   647 => x"a4b05188",
   648 => x"e32d800b",
   649 => x"880c02b8",
   650 => x"050d04a4",
   651 => x"b451909e",
   652 => x"04a4e451",
   653 => x"88e32da5",
   654 => x"9c5188e3",
   655 => x"2da4b051",
   656 => x"88e32da6",
   657 => x"fc08a5dc",
   658 => x"08705471",
   659 => x"87e82953",
   660 => x"5b5699ff",
   661 => x"2d8808a6",
   662 => x"f40c7552",
   663 => x"7987e829",
   664 => x"5199ff2d",
   665 => x"8808a6f8",
   666 => x"0c755279",
   667 => x"84b92951",
   668 => x"99ff2d88",
   669 => x"0880f6ac",
   670 => x"0ca3ac51",
   671 => x"88e32da6",
   672 => x"f40852a3",
   673 => x"dc5188e3",
   674 => x"2da3e451",
   675 => x"88e32da6",
   676 => x"f80852a3",
   677 => x"dc5188e3",
   678 => x"2d80f6ac",
   679 => x"0852a494",
   680 => x"5188e32d",
   681 => x"a4b05188",
   682 => x"e32d800b",
   683 => x"880c02b8",
   684 => x"050d0402",
   685 => x"b805f805",
   686 => x"52805196",
   687 => x"a52d9f53",
   688 => x"a5bc5280",
   689 => x"f688519e",
   690 => x"dd2d7778",
   691 => x"80f5fc0c",
   692 => x"81177081",
   693 => x"ff0680f6",
   694 => x"840b84e0",
   695 => x"2d525856",
   696 => x"5a92e204",
   697 => x"760856b0",
   698 => x"53755276",
   699 => x"519edd2d",
   700 => x"80c10b80",
   701 => x"f6840b84",
   702 => x"e02d5656",
   703 => x"92be04ff",
   704 => x"15707831",
   705 => x"7c0c5980",
   706 => x"59938f04",
   707 => x"02f8050d",
   708 => x"73823270",
   709 => x"09810570",
   710 => x"72078025",
   711 => x"880c5252",
   712 => x"0288050d",
   713 => x"0402f405",
   714 => x"0d747671",
   715 => x"53545271",
   716 => x"822e8338",
   717 => x"83517181",
   718 => x"2e9b3881",
   719 => x"7226a038",
   720 => x"71822ebc",
   721 => x"3871842e",
   722 => x"ac387073",
   723 => x"0c70880c",
   724 => x"028c050d",
   725 => x"0480e40b",
   726 => x"80f5fc08",
   727 => x"258c3880",
   728 => x"730c7088",
   729 => x"0c028c05",
   730 => x"0d048373",
   731 => x"0c70880c",
   732 => x"028c050d",
   733 => x"0482730c",
   734 => x"70880c02",
   735 => x"8c050d04",
   736 => x"81730c70",
   737 => x"880c028c",
   738 => x"050d0402",
   739 => x"fc050d74",
   740 => x"74148205",
   741 => x"710c880c",
   742 => x"0284050d",
   743 => x"0402d805",
   744 => x"0d7b7d7f",
   745 => x"61851270",
   746 => x"822b7511",
   747 => x"70747170",
   748 => x"8405530c",
   749 => x"5a5a5d5b",
   750 => x"760c7980",
   751 => x"f8180c79",
   752 => x"86125257",
   753 => x"585a5a76",
   754 => x"76249938",
   755 => x"76b32982",
   756 => x"2b791151",
   757 => x"53767370",
   758 => x"8405550c",
   759 => x"81145475",
   760 => x"7425f238",
   761 => x"7681cc29",
   762 => x"19fc1108",
   763 => x"8105fc12",
   764 => x"0c7a1970",
   765 => x"089fa013",
   766 => x"0c585685",
   767 => x"0b80f5fc",
   768 => x"0c75880c",
   769 => x"02a8050d",
   770 => x"0402f405",
   771 => x"0d029305",
   772 => x"84e02d51",
   773 => x"80028405",
   774 => x"970584e0",
   775 => x"2d545270",
   776 => x"732e8938",
   777 => x"71880c02",
   778 => x"8c050d04",
   779 => x"7080f680",
   780 => x"0b85802d",
   781 => x"810b880c",
   782 => x"028c050d",
   783 => x"0402dc05",
   784 => x"0d7a7c59",
   785 => x"56820b83",
   786 => x"19555574",
   787 => x"167084e0",
   788 => x"2d7584e0",
   789 => x"2d5b5153",
   790 => x"72792e80",
   791 => x"c73880c1",
   792 => x"0b811681",
   793 => x"16565657",
   794 => x"827525df",
   795 => x"38ffa917",
   796 => x"7081ff06",
   797 => x"55597382",
   798 => x"26833887",
   799 => x"55815376",
   800 => x"80d22e98",
   801 => x"38775275",
   802 => x"519ff62d",
   803 => x"80537288",
   804 => x"08258938",
   805 => x"871580f5",
   806 => x"fc0c8153",
   807 => x"72880c02",
   808 => x"a4050d04",
   809 => x"7280f680",
   810 => x"0b85802d",
   811 => x"827525ff",
   812 => x"9a3898ed",
   813 => x"04940802",
   814 => x"940cfd3d",
   815 => x"0d805394",
   816 => x"088c0508",
   817 => x"52940888",
   818 => x"05085182",
   819 => x"de3f8808",
   820 => x"70880c54",
   821 => x"853d0d94",
   822 => x"0c049408",
   823 => x"02940cfd",
   824 => x"3d0d8153",
   825 => x"94088c05",
   826 => x"08529408",
   827 => x"88050851",
   828 => x"82b93f88",
   829 => x"0870880c",
   830 => x"54853d0d",
   831 => x"940c0494",
   832 => x"0802940c",
   833 => x"f93d0d80",
   834 => x"0b9408fc",
   835 => x"050c9408",
   836 => x"88050880",
   837 => x"25ab3894",
   838 => x"08880508",
   839 => x"30940888",
   840 => x"050c800b",
   841 => x"9408f405",
   842 => x"0c9408fc",
   843 => x"05088838",
   844 => x"810b9408",
   845 => x"f4050c94",
   846 => x"08f40508",
   847 => x"9408fc05",
   848 => x"0c94088c",
   849 => x"05088025",
   850 => x"ab389408",
   851 => x"8c050830",
   852 => x"94088c05",
   853 => x"0c800b94",
   854 => x"08f0050c",
   855 => x"9408fc05",
   856 => x"08883881",
   857 => x"0b9408f0",
   858 => x"050c9408",
   859 => x"f0050894",
   860 => x"08fc050c",
   861 => x"80539408",
   862 => x"8c050852",
   863 => x"94088805",
   864 => x"085181a7",
   865 => x"3f880870",
   866 => x"9408f805",
   867 => x"0c549408",
   868 => x"fc050880",
   869 => x"2e8c3894",
   870 => x"08f80508",
   871 => x"309408f8",
   872 => x"050c9408",
   873 => x"f8050870",
   874 => x"880c5489",
   875 => x"3d0d940c",
   876 => x"04940802",
   877 => x"940cfb3d",
   878 => x"0d800b94",
   879 => x"08fc050c",
   880 => x"94088805",
   881 => x"08802593",
   882 => x"38940888",
   883 => x"05083094",
   884 => x"0888050c",
   885 => x"810b9408",
   886 => x"fc050c94",
   887 => x"088c0508",
   888 => x"80258c38",
   889 => x"94088c05",
   890 => x"08309408",
   891 => x"8c050c81",
   892 => x"5394088c",
   893 => x"05085294",
   894 => x"08880508",
   895 => x"51ad3f88",
   896 => x"08709408",
   897 => x"f8050c54",
   898 => x"9408fc05",
   899 => x"08802e8c",
   900 => x"389408f8",
   901 => x"05083094",
   902 => x"08f8050c",
   903 => x"9408f805",
   904 => x"0870880c",
   905 => x"54873d0d",
   906 => x"940c0494",
   907 => x"0802940c",
   908 => x"fd3d0d81",
   909 => x"0b9408fc",
   910 => x"050c800b",
   911 => x"9408f805",
   912 => x"0c94088c",
   913 => x"05089408",
   914 => x"88050827",
   915 => x"ac389408",
   916 => x"fc050880",
   917 => x"2ea33880",
   918 => x"0b94088c",
   919 => x"05082499",
   920 => x"3894088c",
   921 => x"05081094",
   922 => x"088c050c",
   923 => x"9408fc05",
   924 => x"08109408",
   925 => x"fc050cc9",
   926 => x"399408fc",
   927 => x"0508802e",
   928 => x"80c93894",
   929 => x"088c0508",
   930 => x"94088805",
   931 => x"0826a138",
   932 => x"94088805",
   933 => x"0894088c",
   934 => x"05083194",
   935 => x"0888050c",
   936 => x"9408f805",
   937 => x"089408fc",
   938 => x"05080794",
   939 => x"08f8050c",
   940 => x"9408fc05",
   941 => x"08812a94",
   942 => x"08fc050c",
   943 => x"94088c05",
   944 => x"08812a94",
   945 => x"088c050c",
   946 => x"ffaf3994",
   947 => x"08900508",
   948 => x"802e8f38",
   949 => x"94088805",
   950 => x"08709408",
   951 => x"f4050c51",
   952 => x"8d399408",
   953 => x"f8050870",
   954 => x"9408f405",
   955 => x"0c519408",
   956 => x"f4050888",
   957 => x"0c853d0d",
   958 => x"940c0494",
   959 => x"0802940c",
   960 => x"ff3d0d80",
   961 => x"0b9408fc",
   962 => x"050c9408",
   963 => x"88050881",
   964 => x"06ff1170",
   965 => x"09709408",
   966 => x"8c050806",
   967 => x"9408fc05",
   968 => x"08119408",
   969 => x"fc050c94",
   970 => x"08880508",
   971 => x"812a9408",
   972 => x"88050c94",
   973 => x"088c0508",
   974 => x"1094088c",
   975 => x"050c5151",
   976 => x"51519408",
   977 => x"88050880",
   978 => x"2e8438ff",
   979 => x"bd399408",
   980 => x"fc050870",
   981 => x"880c5183",
   982 => x"3d0d940c",
   983 => x"04fc3d0d",
   984 => x"7670797b",
   985 => x"55555555",
   986 => x"8f72278c",
   987 => x"38727507",
   988 => x"83065170",
   989 => x"802ea738",
   990 => x"ff125271",
   991 => x"ff2e9838",
   992 => x"72708105",
   993 => x"54337470",
   994 => x"81055634",
   995 => x"ff125271",
   996 => x"ff2e0981",
   997 => x"06ea3874",
   998 => x"880c863d",
   999 => x"0d047451",
  1000 => x"72708405",
  1001 => x"54087170",
  1002 => x"8405530c",
  1003 => x"72708405",
  1004 => x"54087170",
  1005 => x"8405530c",
  1006 => x"72708405",
  1007 => x"54087170",
  1008 => x"8405530c",
  1009 => x"72708405",
  1010 => x"54087170",
  1011 => x"8405530c",
  1012 => x"f0125271",
  1013 => x"8f26c938",
  1014 => x"83722795",
  1015 => x"38727084",
  1016 => x"05540871",
  1017 => x"70840553",
  1018 => x"0cfc1252",
  1019 => x"718326ed",
  1020 => x"387054ff",
  1021 => x"8339fb3d",
  1022 => x"0d777970",
  1023 => x"72078306",
  1024 => x"53545270",
  1025 => x"93387173",
  1026 => x"73085456",
  1027 => x"54717308",
  1028 => x"2e80c438",
  1029 => x"73755452",
  1030 => x"71337081",
  1031 => x"ff065254",
  1032 => x"70802e9d",
  1033 => x"38723355",
  1034 => x"70752e09",
  1035 => x"81069538",
  1036 => x"81128114",
  1037 => x"71337081",
  1038 => x"ff065456",
  1039 => x"545270e5",
  1040 => x"38723355",
  1041 => x"7381ff06",
  1042 => x"7581ff06",
  1043 => x"71713188",
  1044 => x"0c525287",
  1045 => x"3d0d0471",
  1046 => x"0970f7fb",
  1047 => x"fdff1406",
  1048 => x"70f88482",
  1049 => x"81800651",
  1050 => x"51517097",
  1051 => x"38841484",
  1052 => x"16710854",
  1053 => x"56547175",
  1054 => x"082edc38",
  1055 => x"73755452",
  1056 => x"ff963980",
  1057 => x"0b880c87",
  1058 => x"3d0d0400",
  1059 => x"00ffffff",
  1060 => x"ff00ffff",
  1061 => x"ffff00ff",
  1062 => x"ffffff00",
  1063 => x"30313233",
  1064 => x"34353637",
  1065 => x"38394142",
  1066 => x"43444546",
  1067 => x"00000000",
  1068 => x"44485259",
  1069 => x"53544f4e",
  1070 => x"45205052",
  1071 => x"4f475241",
  1072 => x"4d2c2053",
  1073 => x"4f4d4520",
  1074 => x"53545249",
  1075 => x"4e470000",
  1076 => x"44485259",
  1077 => x"53544f4e",
  1078 => x"45205052",
  1079 => x"4f475241",
  1080 => x"4d2c2031",
  1081 => x"27535420",
  1082 => x"53545249",
  1083 => x"4e470000",
  1084 => x"44687279",
  1085 => x"73746f6e",
  1086 => x"65204265",
  1087 => x"6e63686d",
  1088 => x"61726b2c",
  1089 => x"20566572",
  1090 => x"73696f6e",
  1091 => x"20322e31",
  1092 => x"20284c61",
  1093 => x"6e677561",
  1094 => x"67653a20",
  1095 => x"43290a00",
  1096 => x"50726f67",
  1097 => x"72616d20",
  1098 => x"636f6d70",
  1099 => x"696c6564",
  1100 => x"20776974",
  1101 => x"68202772",
  1102 => x"65676973",
  1103 => x"74657227",
  1104 => x"20617474",
  1105 => x"72696275",
  1106 => x"74650a00",
  1107 => x"45786563",
  1108 => x"7574696f",
  1109 => x"6e207374",
  1110 => x"61727473",
  1111 => x"2c202564",
  1112 => x"2072756e",
  1113 => x"73207468",
  1114 => x"726f7567",
  1115 => x"68204468",
  1116 => x"72797374",
  1117 => x"6f6e650a",
  1118 => x"00000000",
  1119 => x"44485259",
  1120 => x"53544f4e",
  1121 => x"45205052",
  1122 => x"4f475241",
  1123 => x"4d2c2032",
  1124 => x"274e4420",
  1125 => x"53545249",
  1126 => x"4e470000",
  1127 => x"55736572",
  1128 => x"2074696d",
  1129 => x"653a2025",
  1130 => x"640a0000",
  1131 => x"4d696372",
  1132 => x"6f736563",
  1133 => x"6f6e6473",
  1134 => x"20666f72",
  1135 => x"206f6e65",
  1136 => x"2072756e",
  1137 => x"20746872",
  1138 => x"6f756768",
  1139 => x"20446872",
  1140 => x"7973746f",
  1141 => x"6e653a20",
  1142 => x"00000000",
  1143 => x"2564200a",
  1144 => x"00000000",
  1145 => x"44687279",
  1146 => x"73746f6e",
  1147 => x"65732070",
  1148 => x"65722053",
  1149 => x"65636f6e",
  1150 => x"643a2020",
  1151 => x"20202020",
  1152 => x"20202020",
  1153 => x"20202020",
  1154 => x"20202020",
  1155 => x"20202020",
  1156 => x"00000000",
  1157 => x"56415820",
  1158 => x"4d495053",
  1159 => x"20726174",
  1160 => x"696e6720",
  1161 => x"2a203130",
  1162 => x"3030203d",
  1163 => x"20256420",
  1164 => x"0a000000",
  1165 => x"50726f67",
  1166 => x"72616d20",
  1167 => x"636f6d70",
  1168 => x"696c6564",
  1169 => x"20776974",
  1170 => x"686f7574",
  1171 => x"20277265",
  1172 => x"67697374",
  1173 => x"65722720",
  1174 => x"61747472",
  1175 => x"69627574",
  1176 => x"650a0000",
  1177 => x"4d656173",
  1178 => x"75726564",
  1179 => x"2074696d",
  1180 => x"6520746f",
  1181 => x"6f20736d",
  1182 => x"616c6c20",
  1183 => x"746f206f",
  1184 => x"62746169",
  1185 => x"6e206d65",
  1186 => x"616e696e",
  1187 => x"6766756c",
  1188 => x"20726573",
  1189 => x"756c7473",
  1190 => x"0a000000",
  1191 => x"506c6561",
  1192 => x"73652069",
  1193 => x"6e637265",
  1194 => x"61736520",
  1195 => x"6e756d62",
  1196 => x"6572206f",
  1197 => x"66207275",
  1198 => x"6e730a00",
  1199 => x"44485259",
  1200 => x"53544f4e",
  1201 => x"45205052",
  1202 => x"4f475241",
  1203 => x"4d2c2033",
  1204 => x"27524420",
  1205 => x"53545249",
  1206 => x"4e470000",
  1207 => x"000061a8",
  1208 => x"00000000",
	others => x"00000000"
);

begin

process (clk)
begin
	if (clk'event and clk = '1') then
		if (from_zpu.memAWriteEnable = '1') and (from_zpu.memBWriteEnable = '1') and (from_zpu.memAAddr=from_zpu.memBAddr) and (from_zpu.memAWrite/=from_zpu.memBWrite) then
			report "write collision" severity failure;
		end if;
	
		if (from_zpu.memAWriteEnable = '1') then
			ram(to_integer(unsigned(from_zpu.memAAddr(maxAddrBit downto 2)))) := from_zpu.memAWrite;
			to_zpu.memARead <= from_zpu.memAWrite;
		else
			to_zpu.memARead <= ram(to_integer(unsigned(from_zpu.memAAddr(maxAddrBit downto 2))));
		end if;
	end if;
end process;

process (clk)
begin
	if (clk'event and clk = '1') then
		if (from_zpu.memBWriteEnable = '1') then
			ram(to_integer(unsigned(from_zpu.memBAddr(maxAddrBit downto 2)))) := from_zpu.memBWrite;
			to_zpu.memBRead <= from_zpu.memBWrite;
		else
			to_zpu.memBRead <= ram(to_integer(unsigned(from_zpu.memBAddr(maxAddrBit downto 2))));
		end if;
	end if;
end process;


end arch;

