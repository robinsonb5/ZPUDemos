-- ZPU
--
-- Copyright 2004-2008 oharboe - �yvind Harboe - oyvind.harboe@zylin.com
-- Modified by Alastair M. Robinson for the ZPUFlex project.
--
-- The FreeBSD license
-- 
-- Redistribution and use in source and binary forms, with or without
-- modification, are permitted provided that the following conditions
-- are met:
-- 
-- 1. Redistributions of source code must retain the above copyright
--    notice, this list of conditions and the following disclaimer.
-- 2. Redistributions in binary form must reproduce the above
--    copyright notice, this list of conditions and the following
--    disclaimer in the documentation and/or other materials
--    provided with the distribution.
-- 
-- THIS SOFTWARE IS PROVIDED BY THE ZPU PROJECT ``AS IS'' AND ANY
-- EXPRESS OR IMPLIED WARRANTIES, INCLUDING, BUT NOT LIMITED TO,
-- THE IMPLIED WARRANTIES OF MERCHANTABILITY AND FITNESS FOR A
-- PARTICULAR PURPOSE ARE DISCLAIMED. IN NO EVENT SHALL THE
-- ZPU PROJECT OR CONTRIBUTORS BE LIABLE FOR ANY DIRECT,
-- INDIRECT, INCIDENTAL, SPECIAL, EXEMPLARY, OR CONSEQUENTIAL DAMAGES
-- (INCLUDING, BUT NOT LIMITED TO, PROCUREMENT OF SUBSTITUTE GOODS
-- OR SERVICES; LOSS OF USE, DATA, OR PROFITS; OR BUSINESS INTERRUPTION)
-- HOWEVER CAUSED AND ON ANY THEORY OF LIABILITY, WHETHER IN CONTRACT,
-- STRICT LIABILITY, OR TORT (INCLUDING NEGLIGENCE OR OTHERWISE)
-- ARISING IN ANY WAY OUT OF THE USE OF THIS SOFTWARE, EVEN IF
-- ADVISED OF THE POSSIBILITY OF SUCH DAMAGE.
-- 
-- The views and conclusions contained in the software and documentation
-- are those of the authors and should not be interpreted as representing
-- official policies, either expressed or implied, of the ZPU Project.

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;


library work;
use work.zpupkg.all;

entity Dhrystone_fast_ROM is
generic
	(
		maxAddrBitBRAM : integer := maxAddrBitBRAMLimit -- Specify your actual ROM size to save LEs and unnecessary block RAM usage.
	);
port (
	clk : in std_logic;
	areset : in std_logic := '0';
	from_zpu : in ZPU_ToROM;
	to_zpu : out ZPU_FromROM
);
end Dhrystone_fast_ROM;

architecture arch of Dhrystone_fast_ROM is

type ram_type is array(natural range 0 to ((2**(maxAddrBitBRAM+1))/4)-1) of std_logic_vector(wordSize-1 downto 0);

shared variable ram : ram_type :=
(
     0 => x"0b0b0b88",
     1 => x"e5040000",
     2 => x"00000000",
     3 => x"00000000",
     4 => x"00000000",
     5 => x"00000000",
     6 => x"00000000",
     7 => x"00000000",
     8 => x"88088c08",
     9 => x"90080b0b",
    10 => x"0b88e108",
    11 => x"2d900c8c",
    12 => x"0c880c04",
    13 => x"00000000",
    14 => x"00000000",
    15 => x"00000000",
    16 => x"71fd0608",
    17 => x"72830609",
    18 => x"81058205",
    19 => x"832b2a83",
    20 => x"ffff0652",
    21 => x"04000000",
    22 => x"00000000",
    23 => x"00000000",
    24 => x"71fd0608",
    25 => x"83ffff73",
    26 => x"83060981",
    27 => x"05820583",
    28 => x"2b2b0906",
    29 => x"7383ffff",
    30 => x"0b0b0b0b",
    31 => x"83a50400",
    32 => x"72098105",
    33 => x"72057373",
    34 => x"09060906",
    35 => x"73097306",
    36 => x"070a8106",
    37 => x"53510400",
    38 => x"00000000",
    39 => x"00000000",
    40 => x"72722473",
    41 => x"732e0753",
    42 => x"51040000",
    43 => x"00000000",
    44 => x"00000000",
    45 => x"00000000",
    46 => x"00000000",
    47 => x"00000000",
    48 => x"71737109",
    49 => x"71068106",
    50 => x"09810572",
    51 => x"0a100a72",
    52 => x"0a100a31",
    53 => x"050a8106",
    54 => x"51515351",
    55 => x"04000000",
    56 => x"72722673",
    57 => x"732e0753",
    58 => x"51040000",
    59 => x"00000000",
    60 => x"00000000",
    61 => x"00000000",
    62 => x"00000000",
    63 => x"00000000",
    64 => x"00000000",
    65 => x"00000000",
    66 => x"00000000",
    67 => x"00000000",
    68 => x"00000000",
    69 => x"00000000",
    70 => x"00000000",
    71 => x"00000000",
    72 => x"0b0b0b88",
    73 => x"ba040000",
    74 => x"00000000",
    75 => x"00000000",
    76 => x"00000000",
    77 => x"00000000",
    78 => x"00000000",
    79 => x"00000000",
    80 => x"720a722b",
    81 => x"0a535104",
    82 => x"00000000",
    83 => x"00000000",
    84 => x"00000000",
    85 => x"00000000",
    86 => x"00000000",
    87 => x"00000000",
    88 => x"72729f06",
    89 => x"0981050b",
    90 => x"0b0b889f",
    91 => x"05040000",
    92 => x"00000000",
    93 => x"00000000",
    94 => x"00000000",
    95 => x"00000000",
    96 => x"72722aff",
    97 => x"739f062a",
    98 => x"0974090a",
    99 => x"8106ff05",
   100 => x"06075351",
   101 => x"04000000",
   102 => x"00000000",
   103 => x"00000000",
   104 => x"71715351",
   105 => x"04067383",
   106 => x"06098105",
   107 => x"8205832b",
   108 => x"0b2b0772",
   109 => x"fc060c51",
   110 => x"51040000",
   111 => x"00000000",
   112 => x"72098105",
   113 => x"72050970",
   114 => x"81050906",
   115 => x"0a810653",
   116 => x"51040000",
   117 => x"00000000",
   118 => x"00000000",
   119 => x"00000000",
   120 => x"72098105",
   121 => x"72050970",
   122 => x"81050906",
   123 => x"0a098106",
   124 => x"53510400",
   125 => x"00000000",
   126 => x"00000000",
   127 => x"00000000",
   128 => x"71098105",
   129 => x"52040000",
   130 => x"00000000",
   131 => x"00000000",
   132 => x"00000000",
   133 => x"00000000",
   134 => x"00000000",
   135 => x"00000000",
   136 => x"72720981",
   137 => x"05055351",
   138 => x"04000000",
   139 => x"00000000",
   140 => x"00000000",
   141 => x"00000000",
   142 => x"00000000",
   143 => x"00000000",
   144 => x"72097206",
   145 => x"73730906",
   146 => x"07535104",
   147 => x"00000000",
   148 => x"00000000",
   149 => x"00000000",
   150 => x"00000000",
   151 => x"00000000",
   152 => x"71fc0608",
   153 => x"72830609",
   154 => x"81058305",
   155 => x"1010102a",
   156 => x"81ff0652",
   157 => x"04000000",
   158 => x"00000000",
   159 => x"00000000",
   160 => x"71fc0608",
   161 => x"0b0b0ba2",
   162 => x"c8738306",
   163 => x"10100508",
   164 => x"060b0b0b",
   165 => x"88a20400",
   166 => x"00000000",
   167 => x"00000000",
   168 => x"88088c08",
   169 => x"90087575",
   170 => x"0b0b0b9b",
   171 => x"bb2d5050",
   172 => x"88085690",
   173 => x"0c8c0c88",
   174 => x"0c510400",
   175 => x"00000000",
   176 => x"88088c08",
   177 => x"90087575",
   178 => x"0b0b0b9c",
   179 => x"ed2d5050",
   180 => x"88085690",
   181 => x"0c8c0c88",
   182 => x"0c510400",
   183 => x"00000000",
   184 => x"72097081",
   185 => x"0509060a",
   186 => x"8106ff05",
   187 => x"70547106",
   188 => x"73097274",
   189 => x"05ff0506",
   190 => x"07515151",
   191 => x"04000000",
   192 => x"72097081",
   193 => x"0509060a",
   194 => x"098106ff",
   195 => x"05705471",
   196 => x"06730972",
   197 => x"7405ff05",
   198 => x"06075151",
   199 => x"51040000",
   200 => x"05ff0504",
   201 => x"00000000",
   202 => x"00000000",
   203 => x"00000000",
   204 => x"00000000",
   205 => x"00000000",
   206 => x"00000000",
   207 => x"00000000",
   208 => x"04000000",
   209 => x"00000000",
   210 => x"00000000",
   211 => x"00000000",
   212 => x"00000000",
   213 => x"00000000",
   214 => x"00000000",
   215 => x"00000000",
   216 => x"71810552",
   217 => x"04000000",
   218 => x"00000000",
   219 => x"00000000",
   220 => x"00000000",
   221 => x"00000000",
   222 => x"00000000",
   223 => x"00000000",
   224 => x"04000000",
   225 => x"00000000",
   226 => x"00000000",
   227 => x"00000000",
   228 => x"00000000",
   229 => x"00000000",
   230 => x"00000000",
   231 => x"00000000",
   232 => x"02840572",
   233 => x"10100552",
   234 => x"04000000",
   235 => x"00000000",
   236 => x"00000000",
   237 => x"00000000",
   238 => x"00000000",
   239 => x"00000000",
   240 => x"00000000",
   241 => x"00000000",
   242 => x"00000000",
   243 => x"00000000",
   244 => x"00000000",
   245 => x"00000000",
   246 => x"00000000",
   247 => x"00000000",
   248 => x"717105ff",
   249 => x"05715351",
   250 => x"020d0400",
   251 => x"00000000",
   252 => x"00000000",
   253 => x"00000000",
   254 => x"00000000",
   255 => x"00000000",
   256 => x"10101010",
   257 => x"10101010",
   258 => x"10101010",
   259 => x"10101010",
   260 => x"10101010",
   261 => x"10101010",
   262 => x"10101010",
   263 => x"10101053",
   264 => x"51047381",
   265 => x"ff067383",
   266 => x"06098105",
   267 => x"83051010",
   268 => x"102b0772",
   269 => x"fc060c51",
   270 => x"51047272",
   271 => x"80728106",
   272 => x"ff050972",
   273 => x"06057110",
   274 => x"52720a10",
   275 => x"0a5372ed",
   276 => x"38515153",
   277 => x"51040000",
   278 => x"800488da",
   279 => x"04040000",
   280 => x"00000004",
   281 => x"5da7a070",
   282 => x"80f9e827",
   283 => x"8b388071",
   284 => x"70840553",
   285 => x"0c88e704",
   286 => x"88da5191",
   287 => x"b30402c0",
   288 => x"050d0280",
   289 => x"c4055b80",
   290 => x"707c7084",
   291 => x"055e0872",
   292 => x"5f5f5f58",
   293 => x"7c708405",
   294 => x"5e085780",
   295 => x"5976982a",
   296 => x"77882b58",
   297 => x"5574802e",
   298 => x"848d387b",
   299 => x"802e80c8",
   300 => x"38805c74",
   301 => x"80e42e81",
   302 => x"f9387480",
   303 => x"f82e81f2",
   304 => x"387480e4",
   305 => x"2e81fd38",
   306 => x"7480e426",
   307 => x"80dd3874",
   308 => x"80e32ebb",
   309 => x"38a5518d",
   310 => x"f02d7451",
   311 => x"8df02d82",
   312 => x"18588119",
   313 => x"59837925",
   314 => x"ffb33874",
   315 => x"ffa6387e",
   316 => x"880c0280",
   317 => x"c0050d04",
   318 => x"74a52e09",
   319 => x"81069838",
   320 => x"810b811a",
   321 => x"5a5c8379",
   322 => x"25ff9238",
   323 => x"89eb047a",
   324 => x"841c7108",
   325 => x"575c5674",
   326 => x"518df02d",
   327 => x"8118811a",
   328 => x"5a588379",
   329 => x"25fef638",
   330 => x"89eb0474",
   331 => x"80f32e83",
   332 => x"8f387480",
   333 => x"f82e0981",
   334 => x"06ff9a38",
   335 => x"7d0b0b0b",
   336 => x"a7f00b0b",
   337 => x"0b0ba7a0",
   338 => x"565b5380",
   339 => x"56757e24",
   340 => x"83913872",
   341 => x"81c538b0",
   342 => x"0b0b0b0b",
   343 => x"a7a00b85",
   344 => x"802d8114",
   345 => x"54ff1454",
   346 => x"7384e02d",
   347 => x"7a708105",
   348 => x"5c85802d",
   349 => x"81165673",
   350 => x"0b0b0ba7",
   351 => x"a02e0981",
   352 => x"06e33880",
   353 => x"7a85802d",
   354 => x"750b0b0b",
   355 => x"a7f05753",
   356 => x"ff135480",
   357 => x"7325feca",
   358 => x"38757081",
   359 => x"055784e0",
   360 => x"2d705255",
   361 => x"8df02d81",
   362 => x"1874ff16",
   363 => x"5654588b",
   364 => x"93047a84",
   365 => x"1c710840",
   366 => x"5c537480",
   367 => x"e42e0981",
   368 => x"06fe8538",
   369 => x"7d0b0b0b",
   370 => x"a7f00b0b",
   371 => x"0b0ba7a0",
   372 => x"565b5380",
   373 => x"56757e24",
   374 => x"81fc3872",
   375 => x"818b38b0",
   376 => x"0b0b0b0b",
   377 => x"a7a00b85",
   378 => x"802d8114",
   379 => x"54ff1454",
   380 => x"7384e02d",
   381 => x"7a708105",
   382 => x"5c85802d",
   383 => x"81165673",
   384 => x"0b0b0ba7",
   385 => x"a02e0981",
   386 => x"06e33880",
   387 => x"7a85802d",
   388 => x"750b0b0b",
   389 => x"a7f05753",
   390 => x"8b900490",
   391 => x"5272519c",
   392 => x"ed2d8808",
   393 => x"a2d80584",
   394 => x"e02d7470",
   395 => x"81055685",
   396 => x"802d9052",
   397 => x"72519bbb",
   398 => x"2d880853",
   399 => x"8808dc38",
   400 => x"730b0b0b",
   401 => x"a7a02efe",
   402 => x"ba38ff14",
   403 => x"547384e0",
   404 => x"2d7a7081",
   405 => x"055c8580",
   406 => x"2d811656",
   407 => x"730b0b0b",
   408 => x"a7a02efe",
   409 => x"9e388ae5",
   410 => x"048a5272",
   411 => x"519ced2d",
   412 => x"8808a2d8",
   413 => x"0584e02d",
   414 => x"74708105",
   415 => x"5685802d",
   416 => x"8a527251",
   417 => x"9bbb2d88",
   418 => x"08538808",
   419 => x"dc38730b",
   420 => x"0b0ba7a0",
   421 => x"2efdec38",
   422 => x"ff145473",
   423 => x"84e02d7a",
   424 => x"7081055c",
   425 => x"85802d81",
   426 => x"1656730b",
   427 => x"0b0ba7a0",
   428 => x"2efed838",
   429 => x"8bed0477",
   430 => x"880c0280",
   431 => x"c0050d04",
   432 => x"7a841c71",
   433 => x"08705458",
   434 => x"5c548e91",
   435 => x"2d800bff",
   436 => x"1155538b",
   437 => x"9304ad51",
   438 => x"8df02d7d",
   439 => x"09810553",
   440 => x"8bdb04ad",
   441 => x"518df02d",
   442 => x"7d098105",
   443 => x"538ad304",
   444 => x"02f8050d",
   445 => x"7352c008",
   446 => x"70882a70",
   447 => x"81065151",
   448 => x"5170802e",
   449 => x"f13871c0",
   450 => x"0c71880c",
   451 => x"0288050d",
   452 => x"0402e805",
   453 => x"0d807857",
   454 => x"55757084",
   455 => x"05570853",
   456 => x"80547298",
   457 => x"2a73882b",
   458 => x"54527180",
   459 => x"2ea238c0",
   460 => x"0870882a",
   461 => x"70810651",
   462 => x"51517080",
   463 => x"2ef13871",
   464 => x"c00c8115",
   465 => x"81155555",
   466 => x"837425d6",
   467 => x"3871ca38",
   468 => x"74880c02",
   469 => x"98050d04",
   470 => x"c808880c",
   471 => x"0402fc05",
   472 => x"0d80c10b",
   473 => x"80f7bc0b",
   474 => x"85802d80",
   475 => x"0b80f9d4",
   476 => x"0c70880c",
   477 => x"0284050d",
   478 => x"0402f805",
   479 => x"0d800b80",
   480 => x"f7bc0b84",
   481 => x"e02d5252",
   482 => x"7080c12e",
   483 => x"9d387180",
   484 => x"f9d40807",
   485 => x"80f9d40c",
   486 => x"80c20b80",
   487 => x"f7c00b85",
   488 => x"802d7088",
   489 => x"0c028805",
   490 => x"0d04810b",
   491 => x"80f9d408",
   492 => x"0780f9d4",
   493 => x"0c80c20b",
   494 => x"80f7c00b",
   495 => x"85802d70",
   496 => x"880c0288",
   497 => x"050d0402",
   498 => x"f0050d75",
   499 => x"70088a05",
   500 => x"535380f7",
   501 => x"bc0b84e0",
   502 => x"2d517080",
   503 => x"c12e8c38",
   504 => x"73f03870",
   505 => x"880c0290",
   506 => x"050d04ff",
   507 => x"127080f7",
   508 => x"b8083174",
   509 => x"0c880c02",
   510 => x"90050d04",
   511 => x"02ec050d",
   512 => x"80f7e408",
   513 => x"5574802e",
   514 => x"8c387675",
   515 => x"08710c80",
   516 => x"f7e40856",
   517 => x"548c1553",
   518 => x"80f7b808",
   519 => x"528a5199",
   520 => x"912d7388",
   521 => x"0c029405",
   522 => x"0d0402e8",
   523 => x"050d7770",
   524 => x"085656b0",
   525 => x"5380f7e4",
   526 => x"08527451",
   527 => x"a0992d85",
   528 => x"0b8c170c",
   529 => x"850b8c16",
   530 => x"0c750875",
   531 => x"0c80f7e4",
   532 => x"08547380",
   533 => x"2e8a3873",
   534 => x"08750c80",
   535 => x"f7e40854",
   536 => x"8c145380",
   537 => x"f7b80852",
   538 => x"8a519991",
   539 => x"2d841508",
   540 => x"ae38860b",
   541 => x"8c160c88",
   542 => x"15528816",
   543 => x"085198ab",
   544 => x"2d80f7e4",
   545 => x"08700876",
   546 => x"0c548c15",
   547 => x"7054548a",
   548 => x"52730851",
   549 => x"99912d73",
   550 => x"880c0298",
   551 => x"050d0475",
   552 => x"0854b053",
   553 => x"73527551",
   554 => x"a0992d73",
   555 => x"880c0298",
   556 => x"050d0402",
   557 => x"c8050d80",
   558 => x"f6d00b80",
   559 => x"f7840c80",
   560 => x"f7880b80",
   561 => x"f7e40c80",
   562 => x"f6d00b80",
   563 => x"f7880c80",
   564 => x"0b80f788",
   565 => x"0b84050c",
   566 => x"820b80f7",
   567 => x"880b8805",
   568 => x"0ca80b80",
   569 => x"f7880b8c",
   570 => x"050c9f53",
   571 => x"a2ec5280",
   572 => x"f79851a0",
   573 => x"992d9f53",
   574 => x"a38c5280",
   575 => x"f9b451a0",
   576 => x"992d8a0b",
   577 => x"b59c0ca5",
   578 => x"ec5188fe",
   579 => x"2da3ac51",
   580 => x"88fe2da5",
   581 => x"ec5188fe",
   582 => x"2da79c08",
   583 => x"802e8491",
   584 => x"38a3dc51",
   585 => x"88fe2da5",
   586 => x"ec5188fe",
   587 => x"2da79808",
   588 => x"52a48851",
   589 => x"88fe2dc8",
   590 => x"0870a8bc",
   591 => x"0c568158",
   592 => x"800ba798",
   593 => x"082582dc",
   594 => x"3802ac05",
   595 => x"5b80c10b",
   596 => x"80f7bc0b",
   597 => x"85802d81",
   598 => x"0b80f9d4",
   599 => x"0c80c20b",
   600 => x"80f7c00b",
   601 => x"85802d82",
   602 => x"5c835a9f",
   603 => x"53a4b852",
   604 => x"80f7c451",
   605 => x"a0992d81",
   606 => x"5d800b80",
   607 => x"f7c45380",
   608 => x"f9b45255",
   609 => x"9ac32d88",
   610 => x"08752e09",
   611 => x"81068338",
   612 => x"81557480",
   613 => x"f9d40c7b",
   614 => x"70575574",
   615 => x"8325a138",
   616 => x"74101015",
   617 => x"fd055e02",
   618 => x"b805fc05",
   619 => x"53835275",
   620 => x"5199912d",
   621 => x"811c705d",
   622 => x"70575583",
   623 => x"7524e138",
   624 => x"7d547453",
   625 => x"a8c05280",
   626 => x"f7ec5199",
   627 => x"a32d80f7",
   628 => x"e4087008",
   629 => x"5757b053",
   630 => x"76527551",
   631 => x"a0992d85",
   632 => x"0b8c180c",
   633 => x"850b8c17",
   634 => x"0c760876",
   635 => x"0c80f7e4",
   636 => x"08557480",
   637 => x"2e8a3874",
   638 => x"08760c80",
   639 => x"f7e40855",
   640 => x"8c155380",
   641 => x"f7b80852",
   642 => x"8a519991",
   643 => x"2d841608",
   644 => x"83d83886",
   645 => x"0b8c170c",
   646 => x"88165288",
   647 => x"17085198",
   648 => x"ab2d80f7",
   649 => x"e4087008",
   650 => x"770c578c",
   651 => x"16705455",
   652 => x"8a527408",
   653 => x"5199912d",
   654 => x"80c10b80",
   655 => x"f7c00b84",
   656 => x"e02d5656",
   657 => x"757526a5",
   658 => x"3880c352",
   659 => x"75519a8f",
   660 => x"2d88087d",
   661 => x"2e82e238",
   662 => x"81167081",
   663 => x"ff0680f7",
   664 => x"c00b84e0",
   665 => x"2d525755",
   666 => x"747627dd",
   667 => x"38797c29",
   668 => x"7e53519b",
   669 => x"bb2d8808",
   670 => x"5c88088a",
   671 => x"0580f7bc",
   672 => x"0b84e02d",
   673 => x"80f7b808",
   674 => x"59575575",
   675 => x"80c12e82",
   676 => x"f43878f7",
   677 => x"38811858",
   678 => x"a7980878",
   679 => x"25fdae38",
   680 => x"a8bc0856",
   681 => x"c8087080",
   682 => x"f7800c70",
   683 => x"773170a8",
   684 => x"b80c53a4",
   685 => x"d8525b88",
   686 => x"fe2da8b8",
   687 => x"085680f7",
   688 => x"762580f3",
   689 => x"38a79808",
   690 => x"70537687",
   691 => x"e829525a",
   692 => x"9bbb2d88",
   693 => x"08a8b00c",
   694 => x"75527987",
   695 => x"e829519b",
   696 => x"bb2d8808",
   697 => x"a8b40c75",
   698 => x"527984b9",
   699 => x"29519bbb",
   700 => x"2d880880",
   701 => x"f7e80ca4",
   702 => x"e85188fe",
   703 => x"2da8b008",
   704 => x"52a59851",
   705 => x"88fe2da5",
   706 => x"a05188fe",
   707 => x"2da8b408",
   708 => x"52a59851",
   709 => x"88fe2d80",
   710 => x"f7e80852",
   711 => x"a5d05188",
   712 => x"fe2da5ec",
   713 => x"5188fe2d",
   714 => x"800b880c",
   715 => x"02b8050d",
   716 => x"04a5f051",
   717 => x"92a404a6",
   718 => x"a05188fe",
   719 => x"2da6d851",
   720 => x"88fe2da5",
   721 => x"ec5188fe",
   722 => x"2da8b808",
   723 => x"a7980870",
   724 => x"547187e8",
   725 => x"29535b56",
   726 => x"9bbb2d88",
   727 => x"08a8b00c",
   728 => x"75527987",
   729 => x"e829519b",
   730 => x"bb2d8808",
   731 => x"a8b40c75",
   732 => x"527984b9",
   733 => x"29519bbb",
   734 => x"2d880880",
   735 => x"f7e80ca4",
   736 => x"e85188fe",
   737 => x"2da8b008",
   738 => x"52a59851",
   739 => x"88fe2da5",
   740 => x"a05188fe",
   741 => x"2da8b408",
   742 => x"52a59851",
   743 => x"88fe2d80",
   744 => x"f7e80852",
   745 => x"a5d05188",
   746 => x"fe2da5ec",
   747 => x"5188fe2d",
   748 => x"800b880c",
   749 => x"02b8050d",
   750 => x"0402b805",
   751 => x"f8055280",
   752 => x"5198ab2d",
   753 => x"9f53a6f8",
   754 => x"5280f7c4",
   755 => x"51a0992d",
   756 => x"777880f7",
   757 => x"b80c8117",
   758 => x"7081ff06",
   759 => x"80f7c00b",
   760 => x"84e02d52",
   761 => x"58565a94",
   762 => x"e8047608",
   763 => x"56b05375",
   764 => x"527651a0",
   765 => x"992d80c1",
   766 => x"0b80f7c0",
   767 => x"0b84e02d",
   768 => x"565694c4",
   769 => x"04ff1570",
   770 => x"78317c0c",
   771 => x"59805995",
   772 => x"950402f8",
   773 => x"050d7382",
   774 => x"32700981",
   775 => x"05707207",
   776 => x"8025880c",
   777 => x"52520288",
   778 => x"050d0402",
   779 => x"f4050d74",
   780 => x"76715354",
   781 => x"5271822e",
   782 => x"83388351",
   783 => x"71812e9b",
   784 => x"38817226",
   785 => x"a0387182",
   786 => x"2ebc3871",
   787 => x"842eac38",
   788 => x"70730c70",
   789 => x"880c028c",
   790 => x"050d0480",
   791 => x"e40b80f7",
   792 => x"b808258c",
   793 => x"3880730c",
   794 => x"70880c02",
   795 => x"8c050d04",
   796 => x"83730c70",
   797 => x"880c028c",
   798 => x"050d0482",
   799 => x"730c7088",
   800 => x"0c028c05",
   801 => x"0d048173",
   802 => x"0c70880c",
   803 => x"028c050d",
   804 => x"0402fc05",
   805 => x"0d747414",
   806 => x"8205710c",
   807 => x"880c0284",
   808 => x"050d0402",
   809 => x"d8050d7b",
   810 => x"7d7f6185",
   811 => x"1270822b",
   812 => x"75117074",
   813 => x"71708405",
   814 => x"530c5a5a",
   815 => x"5d5b760c",
   816 => x"7980f818",
   817 => x"0c798612",
   818 => x"5257585a",
   819 => x"5a767624",
   820 => x"993876b3",
   821 => x"29822b79",
   822 => x"11515376",
   823 => x"73708405",
   824 => x"550c8114",
   825 => x"54757425",
   826 => x"f2387681",
   827 => x"cc2919fc",
   828 => x"11088105",
   829 => x"fc120c7a",
   830 => x"1970089f",
   831 => x"a0130c58",
   832 => x"56850b80",
   833 => x"f7b80c75",
   834 => x"880c02a8",
   835 => x"050d0402",
   836 => x"f4050d02",
   837 => x"930584e0",
   838 => x"2d518002",
   839 => x"84059705",
   840 => x"84e02d54",
   841 => x"5270732e",
   842 => x"89387188",
   843 => x"0c028c05",
   844 => x"0d047080",
   845 => x"f7bc0b85",
   846 => x"802d810b",
   847 => x"880c028c",
   848 => x"050d0402",
   849 => x"dc050d7a",
   850 => x"7c595682",
   851 => x"0b831955",
   852 => x"55741670",
   853 => x"84e02d75",
   854 => x"84e02d5b",
   855 => x"51537279",
   856 => x"2e80c738",
   857 => x"80c10b81",
   858 => x"16811656",
   859 => x"56578275",
   860 => x"25df38ff",
   861 => x"a9177081",
   862 => x"ff065559",
   863 => x"73822683",
   864 => x"38875581",
   865 => x"537680d2",
   866 => x"2e983877",
   867 => x"527551a1",
   868 => x"b22d8053",
   869 => x"72880825",
   870 => x"89388715",
   871 => x"80f7b80c",
   872 => x"81537288",
   873 => x"0c02a405",
   874 => x"0d047280",
   875 => x"f7bc0b85",
   876 => x"802d8275",
   877 => x"25ff9a38",
   878 => x"9af30494",
   879 => x"0802940c",
   880 => x"f93d0d80",
   881 => x"0b9408fc",
   882 => x"050c9408",
   883 => x"88050880",
   884 => x"25ab3894",
   885 => x"08880508",
   886 => x"30940888",
   887 => x"050c800b",
   888 => x"9408f405",
   889 => x"0c9408fc",
   890 => x"05088838",
   891 => x"810b9408",
   892 => x"f4050c94",
   893 => x"08f40508",
   894 => x"9408fc05",
   895 => x"0c94088c",
   896 => x"05088025",
   897 => x"ab389408",
   898 => x"8c050830",
   899 => x"94088c05",
   900 => x"0c800b94",
   901 => x"08f0050c",
   902 => x"9408fc05",
   903 => x"08883881",
   904 => x"0b9408f0",
   905 => x"050c9408",
   906 => x"f0050894",
   907 => x"08fc050c",
   908 => x"80539408",
   909 => x"8c050852",
   910 => x"94088805",
   911 => x"085181a7",
   912 => x"3f880870",
   913 => x"9408f805",
   914 => x"0c549408",
   915 => x"fc050880",
   916 => x"2e8c3894",
   917 => x"08f80508",
   918 => x"309408f8",
   919 => x"050c9408",
   920 => x"f8050870",
   921 => x"880c5489",
   922 => x"3d0d940c",
   923 => x"04940802",
   924 => x"940cfb3d",
   925 => x"0d800b94",
   926 => x"08fc050c",
   927 => x"94088805",
   928 => x"08802593",
   929 => x"38940888",
   930 => x"05083094",
   931 => x"0888050c",
   932 => x"810b9408",
   933 => x"fc050c94",
   934 => x"088c0508",
   935 => x"80258c38",
   936 => x"94088c05",
   937 => x"08309408",
   938 => x"8c050c81",
   939 => x"5394088c",
   940 => x"05085294",
   941 => x"08880508",
   942 => x"51ad3f88",
   943 => x"08709408",
   944 => x"f8050c54",
   945 => x"9408fc05",
   946 => x"08802e8c",
   947 => x"389408f8",
   948 => x"05083094",
   949 => x"08f8050c",
   950 => x"9408f805",
   951 => x"0870880c",
   952 => x"54873d0d",
   953 => x"940c0494",
   954 => x"0802940c",
   955 => x"fd3d0d81",
   956 => x"0b9408fc",
   957 => x"050c800b",
   958 => x"9408f805",
   959 => x"0c94088c",
   960 => x"05089408",
   961 => x"88050827",
   962 => x"ac389408",
   963 => x"fc050880",
   964 => x"2ea33880",
   965 => x"0b94088c",
   966 => x"05082499",
   967 => x"3894088c",
   968 => x"05081094",
   969 => x"088c050c",
   970 => x"9408fc05",
   971 => x"08109408",
   972 => x"fc050cc9",
   973 => x"399408fc",
   974 => x"0508802e",
   975 => x"80c93894",
   976 => x"088c0508",
   977 => x"94088805",
   978 => x"0826a138",
   979 => x"94088805",
   980 => x"0894088c",
   981 => x"05083194",
   982 => x"0888050c",
   983 => x"9408f805",
   984 => x"089408fc",
   985 => x"05080794",
   986 => x"08f8050c",
   987 => x"9408fc05",
   988 => x"08812a94",
   989 => x"08fc050c",
   990 => x"94088c05",
   991 => x"08812a94",
   992 => x"088c050c",
   993 => x"ffaf3994",
   994 => x"08900508",
   995 => x"802e8f38",
   996 => x"94088805",
   997 => x"08709408",
   998 => x"f4050c51",
   999 => x"8d399408",
  1000 => x"f8050870",
  1001 => x"9408f405",
  1002 => x"0c519408",
  1003 => x"f4050888",
  1004 => x"0c853d0d",
  1005 => x"940c0494",
  1006 => x"0802940c",
  1007 => x"ff3d0d80",
  1008 => x"0b9408fc",
  1009 => x"050c9408",
  1010 => x"88050881",
  1011 => x"06ff1170",
  1012 => x"09709408",
  1013 => x"8c050806",
  1014 => x"9408fc05",
  1015 => x"08119408",
  1016 => x"fc050c94",
  1017 => x"08880508",
  1018 => x"812a9408",
  1019 => x"88050c94",
  1020 => x"088c0508",
  1021 => x"1094088c",
  1022 => x"050c5151",
  1023 => x"51519408",
  1024 => x"88050880",
  1025 => x"2e8438ff",
  1026 => x"bd399408",
  1027 => x"fc050870",
  1028 => x"880c5183",
  1029 => x"3d0d940c",
  1030 => x"04fc3d0d",
  1031 => x"7670797b",
  1032 => x"55555555",
  1033 => x"8f72278c",
  1034 => x"38727507",
  1035 => x"83065170",
  1036 => x"802ea738",
  1037 => x"ff125271",
  1038 => x"ff2e9838",
  1039 => x"72708105",
  1040 => x"54337470",
  1041 => x"81055634",
  1042 => x"ff125271",
  1043 => x"ff2e0981",
  1044 => x"06ea3874",
  1045 => x"880c863d",
  1046 => x"0d047451",
  1047 => x"72708405",
  1048 => x"54087170",
  1049 => x"8405530c",
  1050 => x"72708405",
  1051 => x"54087170",
  1052 => x"8405530c",
  1053 => x"72708405",
  1054 => x"54087170",
  1055 => x"8405530c",
  1056 => x"72708405",
  1057 => x"54087170",
  1058 => x"8405530c",
  1059 => x"f0125271",
  1060 => x"8f26c938",
  1061 => x"83722795",
  1062 => x"38727084",
  1063 => x"05540871",
  1064 => x"70840553",
  1065 => x"0cfc1252",
  1066 => x"718326ed",
  1067 => x"387054ff",
  1068 => x"8339fb3d",
  1069 => x"0d777970",
  1070 => x"72078306",
  1071 => x"53545270",
  1072 => x"93387173",
  1073 => x"73085456",
  1074 => x"54717308",
  1075 => x"2e80c438",
  1076 => x"73755452",
  1077 => x"71337081",
  1078 => x"ff065254",
  1079 => x"70802e9d",
  1080 => x"38723355",
  1081 => x"70752e09",
  1082 => x"81069538",
  1083 => x"81128114",
  1084 => x"71337081",
  1085 => x"ff065456",
  1086 => x"545270e5",
  1087 => x"38723355",
  1088 => x"7381ff06",
  1089 => x"7581ff06",
  1090 => x"71713188",
  1091 => x"0c525287",
  1092 => x"3d0d0471",
  1093 => x"0970f7fb",
  1094 => x"fdff1406",
  1095 => x"70f88482",
  1096 => x"81800651",
  1097 => x"51517097",
  1098 => x"38841484",
  1099 => x"16710854",
  1100 => x"56547175",
  1101 => x"082edc38",
  1102 => x"73755452",
  1103 => x"ff963980",
  1104 => x"0b880c87",
  1105 => x"3d0d0400",
  1106 => x"00ffffff",
  1107 => x"ff00ffff",
  1108 => x"ffff00ff",
  1109 => x"ffffff00",
  1110 => x"30313233",
  1111 => x"34353637",
  1112 => x"38394142",
  1113 => x"43444546",
  1114 => x"00000000",
  1115 => x"44485259",
  1116 => x"53544f4e",
  1117 => x"45205052",
  1118 => x"4f475241",
  1119 => x"4d2c2053",
  1120 => x"4f4d4520",
  1121 => x"53545249",
  1122 => x"4e470000",
  1123 => x"44485259",
  1124 => x"53544f4e",
  1125 => x"45205052",
  1126 => x"4f475241",
  1127 => x"4d2c2031",
  1128 => x"27535420",
  1129 => x"53545249",
  1130 => x"4e470000",
  1131 => x"44687279",
  1132 => x"73746f6e",
  1133 => x"65204265",
  1134 => x"6e63686d",
  1135 => x"61726b2c",
  1136 => x"20566572",
  1137 => x"73696f6e",
  1138 => x"20322e31",
  1139 => x"20284c61",
  1140 => x"6e677561",
  1141 => x"67653a20",
  1142 => x"43290a00",
  1143 => x"50726f67",
  1144 => x"72616d20",
  1145 => x"636f6d70",
  1146 => x"696c6564",
  1147 => x"20776974",
  1148 => x"68202772",
  1149 => x"65676973",
  1150 => x"74657227",
  1151 => x"20617474",
  1152 => x"72696275",
  1153 => x"74650a00",
  1154 => x"45786563",
  1155 => x"7574696f",
  1156 => x"6e207374",
  1157 => x"61727473",
  1158 => x"2c202564",
  1159 => x"2072756e",
  1160 => x"73207468",
  1161 => x"726f7567",
  1162 => x"68204468",
  1163 => x"72797374",
  1164 => x"6f6e650a",
  1165 => x"00000000",
  1166 => x"44485259",
  1167 => x"53544f4e",
  1168 => x"45205052",
  1169 => x"4f475241",
  1170 => x"4d2c2032",
  1171 => x"274e4420",
  1172 => x"53545249",
  1173 => x"4e470000",
  1174 => x"55736572",
  1175 => x"2074696d",
  1176 => x"653a2025",
  1177 => x"640a0000",
  1178 => x"4d696372",
  1179 => x"6f736563",
  1180 => x"6f6e6473",
  1181 => x"20666f72",
  1182 => x"206f6e65",
  1183 => x"2072756e",
  1184 => x"20746872",
  1185 => x"6f756768",
  1186 => x"20446872",
  1187 => x"7973746f",
  1188 => x"6e653a20",
  1189 => x"00000000",
  1190 => x"2564200a",
  1191 => x"00000000",
  1192 => x"44687279",
  1193 => x"73746f6e",
  1194 => x"65732070",
  1195 => x"65722053",
  1196 => x"65636f6e",
  1197 => x"643a2020",
  1198 => x"20202020",
  1199 => x"20202020",
  1200 => x"20202020",
  1201 => x"20202020",
  1202 => x"20202020",
  1203 => x"00000000",
  1204 => x"56415820",
  1205 => x"4d495053",
  1206 => x"20726174",
  1207 => x"696e6720",
  1208 => x"2a203130",
  1209 => x"3030203d",
  1210 => x"20256420",
  1211 => x"0a000000",
  1212 => x"50726f67",
  1213 => x"72616d20",
  1214 => x"636f6d70",
  1215 => x"696c6564",
  1216 => x"20776974",
  1217 => x"686f7574",
  1218 => x"20277265",
  1219 => x"67697374",
  1220 => x"65722720",
  1221 => x"61747472",
  1222 => x"69627574",
  1223 => x"650a0000",
  1224 => x"4d656173",
  1225 => x"75726564",
  1226 => x"2074696d",
  1227 => x"6520746f",
  1228 => x"6f20736d",
  1229 => x"616c6c20",
  1230 => x"746f206f",
  1231 => x"62746169",
  1232 => x"6e206d65",
  1233 => x"616e696e",
  1234 => x"6766756c",
  1235 => x"20726573",
  1236 => x"756c7473",
  1237 => x"0a000000",
  1238 => x"506c6561",
  1239 => x"73652069",
  1240 => x"6e637265",
  1241 => x"61736520",
  1242 => x"6e756d62",
  1243 => x"6572206f",
  1244 => x"66207275",
  1245 => x"6e730a00",
  1246 => x"44485259",
  1247 => x"53544f4e",
  1248 => x"45205052",
  1249 => x"4f475241",
  1250 => x"4d2c2033",
  1251 => x"27524420",
  1252 => x"53545249",
  1253 => x"4e470000",
  1254 => x"000061a8",
  1255 => x"00000000",
	others => x"00000000"
);

begin

process (clk)
begin
	if (clk'event and clk = '1') then
		if (from_zpu.memAWriteEnable = '1') and (from_zpu.memBWriteEnable = '1') and (from_zpu.memAAddr=from_zpu.memBAddr) and (from_zpu.memAWrite/=from_zpu.memBWrite) then
			report "write collision" severity failure;
		end if;
	
		if (from_zpu.memAWriteEnable = '1') then
			ram(to_integer(unsigned(from_zpu.memAAddr(maxAddrBitBRAM downto 2)))) := from_zpu.memAWrite;
			to_zpu.memARead <= from_zpu.memAWrite;
		else
			to_zpu.memARead <= ram(to_integer(unsigned(from_zpu.memAAddr(maxAddrBitBRAM downto 2))));
		end if;
	end if;
end process;

process (clk)
begin
	if (clk'event and clk = '1') then
		if (from_zpu.memBWriteEnable = '1') then
			ram(to_integer(unsigned(from_zpu.memBAddr(maxAddrBitBRAM downto 2)))) := from_zpu.memBWrite;
			to_zpu.memBRead <= from_zpu.memBWrite;
		else
			to_zpu.memBRead <= ram(to_integer(unsigned(from_zpu.memBAddr(maxAddrBitBRAM downto 2))));
		end if;
	end if;
end process;


end arch;

