-- ZPU
--
-- Copyright 2004-2008 oharboe - �yvind Harboe - oyvind.harboe@zylin.com
-- Modified by Alastair M. Robinson for the ZPUFlex project.
--
-- The FreeBSD license
-- 
-- Redistribution and use in source and binary forms, with or without
-- modification, are permitted provided that the following conditions
-- are met:
-- 
-- 1. Redistributions of source code must retain the above copyright
--    notice, this list of conditions and the following disclaimer.
-- 2. Redistributions in binary form must reproduce the above
--    copyright notice, this list of conditions and the following
--    disclaimer in the documentation and/or other materials
--    provided with the distribution.
-- 
-- THIS SOFTWARE IS PROVIDED BY THE ZPU PROJECT ``AS IS'' AND ANY
-- EXPRESS OR IMPLIED WARRANTIES, INCLUDING, BUT NOT LIMITED TO,
-- THE IMPLIED WARRANTIES OF MERCHANTABILITY AND FITNESS FOR A
-- PARTICULAR PURPOSE ARE DISCLAIMED. IN NO EVENT SHALL THE
-- ZPU PROJECT OR CONTRIBUTORS BE LIABLE FOR ANY DIRECT,
-- INDIRECT, INCIDENTAL, SPECIAL, EXEMPLARY, OR CONSEQUENTIAL DAMAGES
-- (INCLUDING, BUT NOT LIMITED TO, PROCUREMENT OF SUBSTITUTE GOODS
-- OR SERVICES; LOSS OF USE, DATA, OR PROFITS; OR BUSINESS INTERRUPTION)
-- HOWEVER CAUSED AND ON ANY THEORY OF LIABILITY, WHETHER IN CONTRACT,
-- STRICT LIABILITY, OR TORT (INCLUDING NEGLIGENCE OR OTHERWISE)
-- ARISING IN ANY WAY OUT OF THE USE OF THIS SOFTWARE, EVEN IF
-- ADVISED OF THE POSSIBILITY OF SUCH DAMAGE.
-- 
-- The views and conclusions contained in the software and documentation
-- are those of the authors and should not be interpreted as representing
-- official policies, either expressed or implied, of the ZPU Project.

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;


library work;
use work.zpu_config.all;
use work.zpupkg.all;

entity Interrupt_ROM is
generic
	(
		maxAddrBitBRAM : integer := maxAddrBitBRAMLimit -- Specify your actual ROM size to save LEs and unnecessary block RAM usage.
	);
port (
	clk : in std_logic;
	areset : in std_logic := '0';
	from_zpu : in ZPU_ToROM;
	to_zpu : out ZPU_FromROM
);
end Interrupt_ROM;

architecture arch of Interrupt_ROM is

type ram_type is array(natural range 0 to ((2**(maxAddrBitBRAM+1))/4)-1) of std_logic_vector(wordSize-1 downto 0);

shared variable ram : ram_type :=
(
     0 => x"0b0b0b88",
     1 => x"e5040000",
     2 => x"00000000",
     3 => x"00000000",
     4 => x"00000000",
     5 => x"00000000",
     6 => x"00000000",
     7 => x"00000000",
     8 => x"88088c08",
     9 => x"90080b0b",
    10 => x"0b88e108",
    11 => x"2d900c8c",
    12 => x"0c880c04",
    13 => x"00000000",
    14 => x"00000000",
    15 => x"00000000",
    16 => x"71fd0608",
    17 => x"72830609",
    18 => x"81058205",
    19 => x"832b2a83",
    20 => x"ffff0652",
    21 => x"04000000",
    22 => x"00000000",
    23 => x"00000000",
    24 => x"71fd0608",
    25 => x"83ffff73",
    26 => x"83060981",
    27 => x"05820583",
    28 => x"2b2b0906",
    29 => x"7383ffff",
    30 => x"0b0b0b0b",
    31 => x"83a50400",
    32 => x"72098105",
    33 => x"72057373",
    34 => x"09060906",
    35 => x"73097306",
    36 => x"070a8106",
    37 => x"53510400",
    38 => x"00000000",
    39 => x"00000000",
    40 => x"72722473",
    41 => x"732e0753",
    42 => x"51040000",
    43 => x"00000000",
    44 => x"00000000",
    45 => x"00000000",
    46 => x"00000000",
    47 => x"00000000",
    48 => x"71737109",
    49 => x"71068106",
    50 => x"09810572",
    51 => x"0a100a72",
    52 => x"0a100a31",
    53 => x"050a8106",
    54 => x"51515351",
    55 => x"04000000",
    56 => x"72722673",
    57 => x"732e0753",
    58 => x"51040000",
    59 => x"00000000",
    60 => x"00000000",
    61 => x"00000000",
    62 => x"00000000",
    63 => x"00000000",
    64 => x"00000000",
    65 => x"00000000",
    66 => x"00000000",
    67 => x"00000000",
    68 => x"00000000",
    69 => x"00000000",
    70 => x"00000000",
    71 => x"00000000",
    72 => x"0b0b0b88",
    73 => x"ba040000",
    74 => x"00000000",
    75 => x"00000000",
    76 => x"00000000",
    77 => x"00000000",
    78 => x"00000000",
    79 => x"00000000",
    80 => x"720a722b",
    81 => x"0a535104",
    82 => x"00000000",
    83 => x"00000000",
    84 => x"00000000",
    85 => x"00000000",
    86 => x"00000000",
    87 => x"00000000",
    88 => x"72729f06",
    89 => x"0981050b",
    90 => x"0b0b889f",
    91 => x"05040000",
    92 => x"00000000",
    93 => x"00000000",
    94 => x"00000000",
    95 => x"00000000",
    96 => x"72722aff",
    97 => x"739f062a",
    98 => x"0974090a",
    99 => x"8106ff05",
   100 => x"06075351",
   101 => x"04000000",
   102 => x"00000000",
   103 => x"00000000",
   104 => x"71715351",
   105 => x"04067383",
   106 => x"06098105",
   107 => x"8205832b",
   108 => x"0b2b0772",
   109 => x"fc060c51",
   110 => x"51040000",
   111 => x"00000000",
   112 => x"72098105",
   113 => x"72050970",
   114 => x"81050906",
   115 => x"0a810653",
   116 => x"51040000",
   117 => x"00000000",
   118 => x"00000000",
   119 => x"00000000",
   120 => x"72098105",
   121 => x"72050970",
   122 => x"81050906",
   123 => x"0a098106",
   124 => x"53510400",
   125 => x"00000000",
   126 => x"00000000",
   127 => x"00000000",
   128 => x"71098105",
   129 => x"52040000",
   130 => x"00000000",
   131 => x"00000000",
   132 => x"00000000",
   133 => x"00000000",
   134 => x"00000000",
   135 => x"00000000",
   136 => x"72720981",
   137 => x"05055351",
   138 => x"04000000",
   139 => x"00000000",
   140 => x"00000000",
   141 => x"00000000",
   142 => x"00000000",
   143 => x"00000000",
   144 => x"72097206",
   145 => x"73730906",
   146 => x"07535104",
   147 => x"00000000",
   148 => x"00000000",
   149 => x"00000000",
   150 => x"00000000",
   151 => x"00000000",
   152 => x"71fc0608",
   153 => x"72830609",
   154 => x"81058305",
   155 => x"1010102a",
   156 => x"81ff0652",
   157 => x"04000000",
   158 => x"00000000",
   159 => x"00000000",
   160 => x"71fc0608",
   161 => x"0b0b0b90",
   162 => x"ec738306",
   163 => x"10100508",
   164 => x"060b0b0b",
   165 => x"88a20400",
   166 => x"00000000",
   167 => x"00000000",
   168 => x"88088c08",
   169 => x"90087575",
   170 => x"0b0b0b8c",
   171 => x"f02d5050",
   172 => x"88085690",
   173 => x"0c8c0c88",
   174 => x"0c510400",
   175 => x"00000000",
   176 => x"88088c08",
   177 => x"90087575",
   178 => x"0b0b0b8e",
   179 => x"a22d5050",
   180 => x"88085690",
   181 => x"0c8c0c88",
   182 => x"0c510400",
   183 => x"00000000",
   184 => x"72097081",
   185 => x"0509060a",
   186 => x"8106ff05",
   187 => x"70547106",
   188 => x"73097274",
   189 => x"05ff0506",
   190 => x"07515151",
   191 => x"04000000",
   192 => x"72097081",
   193 => x"0509060a",
   194 => x"098106ff",
   195 => x"05705471",
   196 => x"06730972",
   197 => x"7405ff05",
   198 => x"06075151",
   199 => x"51040000",
   200 => x"05ff0504",
   201 => x"00000000",
   202 => x"00000000",
   203 => x"00000000",
   204 => x"00000000",
   205 => x"00000000",
   206 => x"00000000",
   207 => x"00000000",
   208 => x"04000000",
   209 => x"00000000",
   210 => x"00000000",
   211 => x"00000000",
   212 => x"00000000",
   213 => x"00000000",
   214 => x"00000000",
   215 => x"00000000",
   216 => x"71810552",
   217 => x"04000000",
   218 => x"00000000",
   219 => x"00000000",
   220 => x"00000000",
   221 => x"00000000",
   222 => x"00000000",
   223 => x"00000000",
   224 => x"00000000",
   225 => x"00000000",
   226 => x"00000000",
   227 => x"00000000",
   228 => x"00000000",
   229 => x"00000000",
   230 => x"00000000",
   231 => x"00000000",
   232 => x"02840572",
   233 => x"10100552",
   234 => x"04000000",
   235 => x"00000000",
   236 => x"00000000",
   237 => x"00000000",
   238 => x"00000000",
   239 => x"00000000",
   240 => x"00000000",
   241 => x"00000000",
   242 => x"00000000",
   243 => x"00000000",
   244 => x"00000000",
   245 => x"00000000",
   246 => x"00000000",
   247 => x"00000000",
   248 => x"717105ff",
   249 => x"05715351",
   250 => x"020d0400",
   251 => x"00000000",
   252 => x"00000000",
   253 => x"00000000",
   254 => x"00000000",
   255 => x"00000000",
   256 => x"10101010",
   257 => x"10101010",
   258 => x"10101010",
   259 => x"10101010",
   260 => x"10101010",
   261 => x"10101010",
   262 => x"10101010",
   263 => x"10101053",
   264 => x"51047381",
   265 => x"ff067383",
   266 => x"06098105",
   267 => x"83051010",
   268 => x"102b0772",
   269 => x"fc060c51",
   270 => x"51047272",
   271 => x"80728106",
   272 => x"ff050972",
   273 => x"06057110",
   274 => x"52720a10",
   275 => x"0a5372ed",
   276 => x"38515153",
   277 => x"51040000",
   278 => x"800488da",
   279 => x"04040000",
   280 => x"00000004",
   281 => x"5d88da0b",
   282 => x"8cba04f0",
   283 => x"3d0d933d",
   284 => x"0b0b0b92",
   285 => x"bc5d5780",
   286 => x"77708405",
   287 => x"59087140",
   288 => x"40597e70",
   289 => x"84054008",
   290 => x"5b805d7a",
   291 => x"982a7b88",
   292 => x"2b5c5675",
   293 => x"86387840",
   294 => x"81f7397d",
   295 => x"802e81d1",
   296 => x"38805e75",
   297 => x"80e42e9b",
   298 => x"387580e4",
   299 => x"268b3875",
   300 => x"80e32e81",
   301 => x"89388190",
   302 => x"397580f3",
   303 => x"2e80ee38",
   304 => x"81863976",
   305 => x"84187108",
   306 => x"0b0b0b92",
   307 => x"bc0b0b0b",
   308 => x"0b91ec62",
   309 => x"5d595d56",
   310 => x"58537380",
   311 => x"258938ad",
   312 => x"5181b53f",
   313 => x"73305473",
   314 => x"8e38b00b",
   315 => x"0b0b0b91",
   316 => x"ec348115",
   317 => x"55a0398a",
   318 => x"743690fc",
   319 => x"05537233",
   320 => x"75708105",
   321 => x"57348a74",
   322 => x"355473eb",
   323 => x"38740b0b",
   324 => x"0b91ec2e",
   325 => x"9138ff15",
   326 => x"5574337a",
   327 => x"7081055c",
   328 => x"34811858",
   329 => x"e839807a",
   330 => x"347754ab",
   331 => x"39768418",
   332 => x"71087054",
   333 => x"5e585380",
   334 => x"fe3f7d54",
   335 => x"9a397684",
   336 => x"18710858",
   337 => x"5853b639",
   338 => x"a55180cc",
   339 => x"3f755180",
   340 => x"c73f8219",
   341 => x"59ae3973",
   342 => x"ff155553",
   343 => x"807325a4",
   344 => x"387b7081",
   345 => x"055d3370",
   346 => x"5256ad3f",
   347 => x"811959e7",
   348 => x"3975a52e",
   349 => x"09810685",
   350 => x"38815e88",
   351 => x"39755198",
   352 => x"3f811959",
   353 => x"811d5d83",
   354 => x"7d25fdff",
   355 => x"3875fdf2",
   356 => x"387f880c",
   357 => x"923d0d04",
   358 => x"ff3d0d73",
   359 => x"52c00870",
   360 => x"882a7081",
   361 => x"06515151",
   362 => x"70802ef1",
   363 => x"3871c00c",
   364 => x"71880c83",
   365 => x"3d0d04fb",
   366 => x"3d0d8078",
   367 => x"57557570",
   368 => x"84055708",
   369 => x"53805472",
   370 => x"982a7388",
   371 => x"2b545271",
   372 => x"802ea238",
   373 => x"c0087088",
   374 => x"2a708106",
   375 => x"51515170",
   376 => x"802ef138",
   377 => x"71c00c81",
   378 => x"15811555",
   379 => x"55837425",
   380 => x"d63871ca",
   381 => x"3874880c",
   382 => x"873d0d04",
   383 => x"7188e10c",
   384 => x"04ffb008",
   385 => x"880c0481",
   386 => x"0bffb00c",
   387 => x"04800bff",
   388 => x"b00c04ff",
   389 => x"3d0df63f",
   390 => x"e83f92fc",
   391 => x"08813270",
   392 => x"92fc0c52",
   393 => x"71802e86",
   394 => x"38919051",
   395 => x"8439919c",
   396 => x"51ff843f",
   397 => x"d23f833d",
   398 => x"0d04803d",
   399 => x"0d800b92",
   400 => x"fc0c91a8",
   401 => x"51fef03f",
   402 => x"800bf884",
   403 => x"0c868da0",
   404 => x"0bf8880c",
   405 => x"91c051fe",
   406 => x"de3f8c93",
   407 => x"51ff9d3f",
   408 => x"ffa53f91",
   409 => x"d851fecf",
   410 => x"3f810bf8",
   411 => x"800cff39",
   412 => x"94080294",
   413 => x"0cf93d0d",
   414 => x"800b9408",
   415 => x"fc050c94",
   416 => x"08880508",
   417 => x"8025ab38",
   418 => x"94088805",
   419 => x"08309408",
   420 => x"88050c80",
   421 => x"0b9408f4",
   422 => x"050c9408",
   423 => x"fc050888",
   424 => x"38810b94",
   425 => x"08f4050c",
   426 => x"9408f405",
   427 => x"089408fc",
   428 => x"050c9408",
   429 => x"8c050880",
   430 => x"25ab3894",
   431 => x"088c0508",
   432 => x"3094088c",
   433 => x"050c800b",
   434 => x"9408f005",
   435 => x"0c9408fc",
   436 => x"05088838",
   437 => x"810b9408",
   438 => x"f0050c94",
   439 => x"08f00508",
   440 => x"9408fc05",
   441 => x"0c805394",
   442 => x"088c0508",
   443 => x"52940888",
   444 => x"05085181",
   445 => x"a73f8808",
   446 => x"709408f8",
   447 => x"050c5494",
   448 => x"08fc0508",
   449 => x"802e8c38",
   450 => x"9408f805",
   451 => x"08309408",
   452 => x"f8050c94",
   453 => x"08f80508",
   454 => x"70880c54",
   455 => x"893d0d94",
   456 => x"0c049408",
   457 => x"02940cfb",
   458 => x"3d0d800b",
   459 => x"9408fc05",
   460 => x"0c940888",
   461 => x"05088025",
   462 => x"93389408",
   463 => x"88050830",
   464 => x"94088805",
   465 => x"0c810b94",
   466 => x"08fc050c",
   467 => x"94088c05",
   468 => x"0880258c",
   469 => x"3894088c",
   470 => x"05083094",
   471 => x"088c050c",
   472 => x"81539408",
   473 => x"8c050852",
   474 => x"94088805",
   475 => x"0851ad3f",
   476 => x"88087094",
   477 => x"08f8050c",
   478 => x"549408fc",
   479 => x"0508802e",
   480 => x"8c389408",
   481 => x"f8050830",
   482 => x"9408f805",
   483 => x"0c9408f8",
   484 => x"05087088",
   485 => x"0c54873d",
   486 => x"0d940c04",
   487 => x"94080294",
   488 => x"0cfd3d0d",
   489 => x"810b9408",
   490 => x"fc050c80",
   491 => x"0b9408f8",
   492 => x"050c9408",
   493 => x"8c050894",
   494 => x"08880508",
   495 => x"27ac3894",
   496 => x"08fc0508",
   497 => x"802ea338",
   498 => x"800b9408",
   499 => x"8c050824",
   500 => x"99389408",
   501 => x"8c050810",
   502 => x"94088c05",
   503 => x"0c9408fc",
   504 => x"05081094",
   505 => x"08fc050c",
   506 => x"c9399408",
   507 => x"fc050880",
   508 => x"2e80c938",
   509 => x"94088c05",
   510 => x"08940888",
   511 => x"050826a1",
   512 => x"38940888",
   513 => x"05089408",
   514 => x"8c050831",
   515 => x"94088805",
   516 => x"0c9408f8",
   517 => x"05089408",
   518 => x"fc050807",
   519 => x"9408f805",
   520 => x"0c9408fc",
   521 => x"0508812a",
   522 => x"9408fc05",
   523 => x"0c94088c",
   524 => x"0508812a",
   525 => x"94088c05",
   526 => x"0cffaf39",
   527 => x"94089005",
   528 => x"08802e8f",
   529 => x"38940888",
   530 => x"05087094",
   531 => x"08f4050c",
   532 => x"518d3994",
   533 => x"08f80508",
   534 => x"709408f4",
   535 => x"050c5194",
   536 => x"08f40508",
   537 => x"880c853d",
   538 => x"0d940c04",
   539 => x"00ffffff",
   540 => x"ff00ffff",
   541 => x"ffff00ff",
   542 => x"ffffff00",
   543 => x"30313233",
   544 => x"34353637",
   545 => x"38394142",
   546 => x"43444546",
   547 => x"00000000",
   548 => x"5469636b",
   549 => x"2e2e2e0a",
   550 => x"00000000",
   551 => x"546f636b",
   552 => x"2e2e2e0a",
   553 => x"00000000",
   554 => x"53657474",
   555 => x"696e6720",
   556 => x"75702074",
   557 => x"696d6572",
   558 => x"2e2e2e0a",
   559 => x"00000000",
   560 => x"456e6162",
   561 => x"6c696e67",
   562 => x"20696e74",
   563 => x"65727275",
   564 => x"7074732e",
   565 => x"2e2e0a00",
   566 => x"456e6162",
   567 => x"6c696e67",
   568 => x"2074696d",
   569 => x"65722e2e",
   570 => x"2e0a002e",
	others => x"00000000"
);

begin

process (clk)
begin
	if (clk'event and clk = '1') then
		if (from_zpu.memAWriteEnable = '1') and (from_zpu.memBWriteEnable = '1') and (from_zpu.memAAddr=from_zpu.memBAddr) and (from_zpu.memAWrite/=from_zpu.memBWrite) then
			report "write collision" severity failure;
		end if;
	
		if (from_zpu.memAWriteEnable = '1') then
			ram(to_integer(unsigned(from_zpu.memAAddr(maxAddrBitBRAM downto 2)))) := from_zpu.memAWrite;
			to_zpu.memARead <= from_zpu.memAWrite;
		else
			to_zpu.memARead <= ram(to_integer(unsigned(from_zpu.memAAddr(maxAddrBitBRAM downto 2))));
		end if;
	end if;
end process;

process (clk)
begin
	if (clk'event and clk = '1') then
		if (from_zpu.memBWriteEnable = '1') then
			ram(to_integer(unsigned(from_zpu.memBAddr(maxAddrBitBRAM downto 2)))) := from_zpu.memBWrite;
			to_zpu.memBRead <= from_zpu.memBWrite;
		else
			to_zpu.memBRead <= ram(to_integer(unsigned(from_zpu.memBAddr(maxAddrBitBRAM downto 2))));
		end if;
	end if;
end process;


end arch;

