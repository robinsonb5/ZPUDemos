-- ZPU
--
-- Copyright 2004-2008 oharboe - �yvind Harboe - oyvind.harboe@zylin.com
-- Modified by Alastair M. Robinson for the ZPUFlex project.
--
-- The FreeBSD license
-- 
-- Redistribution and use in source and binary forms, with or without
-- modification, are permitted provided that the following conditions
-- are met:
-- 
-- 1. Redistributions of source code must retain the above copyright
--    notice, this list of conditions and the following disclaimer.
-- 2. Redistributions in binary form must reproduce the above
--    copyright notice, this list of conditions and the following
--    disclaimer in the documentation and/or other materials
--    provided with the distribution.
-- 
-- THIS SOFTWARE IS PROVIDED BY THE ZPU PROJECT ``AS IS'' AND ANY
-- EXPRESS OR IMPLIED WARRANTIES, INCLUDING, BUT NOT LIMITED TO,
-- THE IMPLIED WARRANTIES OF MERCHANTABILITY AND FITNESS FOR A
-- PARTICULAR PURPOSE ARE DISCLAIMED. IN NO EVENT SHALL THE
-- ZPU PROJECT OR CONTRIBUTORS BE LIABLE FOR ANY DIRECT,
-- INDIRECT, INCIDENTAL, SPECIAL, EXEMPLARY, OR CONSEQUENTIAL DAMAGES
-- (INCLUDING, BUT NOT LIMITED TO, PROCUREMENT OF SUBSTITUTE GOODS
-- OR SERVICES; LOSS OF USE, DATA, OR PROFITS; OR BUSINESS INTERRUPTION)
-- HOWEVER CAUSED AND ON ANY THEORY OF LIABILITY, WHETHER IN CONTRACT,
-- STRICT LIABILITY, OR TORT (INCLUDING NEGLIGENCE OR OTHERWISE)
-- ARISING IN ANY WAY OUT OF THE USE OF THIS SOFTWARE, EVEN IF
-- ADVISED OF THE POSSIBILITY OF SUCH DAMAGE.
-- 
-- The views and conclusions contained in the software and documentation
-- are those of the authors and should not be interpreted as representing
-- official policies, either expressed or implied, of the ZPU Project.

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;


library work;
use work.zpu_config.all;
use work.zpupkg.all;

entity SDRAMTest_ROM is
generic
	(
		maxAddrBit : integer := maxAddrBitBRAMLimit -- Specify your actual ROM size to save LEs and unnecessary block RAM usage.
	);
port (
	clk : in std_logic;
	areset : in std_logic := '0';
	from_zpu : in ZPU_ToROM;
	to_zpu : out ZPU_FromROM
);
end SDRAMTest_ROM;

architecture arch of SDRAMTest_ROM is

type ram_type is array(natural range 0 to ((2**(maxAddrBit+1))/4)-1) of std_logic_vector(wordSize-1 downto 0);

shared variable ram : ram_type :=
(
     0 => x"0ba08080",
     1 => x"e2040000",
     2 => x"8004a080",
     3 => x"808a0471",
     4 => x"fd060872",
     5 => x"83060981",
     6 => x"05820583",
     7 => x"2b2a83ff",
     8 => x"ff065204",
     9 => x"71fc0608",
    10 => x"72830609",
    11 => x"81058305",
    12 => x"1010102a",
    13 => x"81ff0652",
    14 => x"0471fc06",
    15 => x"080ba080",
    16 => x"8ee87383",
    17 => x"06101005",
    18 => x"08067381",
    19 => x"ff067383",
    20 => x"06098105",
    21 => x"83051010",
    22 => x"102b0772",
    23 => x"fc060c51",
    24 => x"5104a080",
    25 => x"808a0ba0",
    26 => x"808be804",
    27 => x"0002c005",
    28 => x"0d0280c4",
    29 => x"05a08095",
    30 => x"d45c5c80",
    31 => x"7c708405",
    32 => x"5e08715f",
    33 => x"5f587d70",
    34 => x"84055f08",
    35 => x"57805a76",
    36 => x"982a7788",
    37 => x"2b585574",
    38 => x"802e8295",
    39 => x"387c802e",
    40 => x"80c23880",
    41 => x"5d7480e4",
    42 => x"2e81b638",
    43 => x"7480e426",
    44 => x"80eb3874",
    45 => x"80e32e80",
    46 => x"c438a551",
    47 => x"a08083bd",
    48 => x"2d7451a0",
    49 => x"8083bd2d",
    50 => x"82185881",
    51 => x"1a5a837a",
    52 => x"25ffbc38",
    53 => x"74ffaf38",
    54 => x"7ea08094",
    55 => x"f40c0280",
    56 => x"c0050d04",
    57 => x"74a52e09",
    58 => x"81069a38",
    59 => x"810b811b",
    60 => x"5b5d837a",
    61 => x"25ff9838",
    62 => x"a08081d4",
    63 => x"047b841d",
    64 => x"7108575d",
    65 => x"547451a0",
    66 => x"8083bd2d",
    67 => x"8118811b",
    68 => x"5b58837a",
    69 => x"25fef838",
    70 => x"a08081d4",
    71 => x"047480f3",
    72 => x"2e098106",
    73 => x"ff94387b",
    74 => x"841d7108",
    75 => x"70545d5d",
    76 => x"53a08083",
    77 => x"e12d800b",
    78 => x"ff115452",
    79 => x"807225ff",
    80 => x"8a387a70",
    81 => x"81055ca0",
    82 => x"8080a42d",
    83 => x"705255a0",
    84 => x"8083bd2d",
    85 => x"811873ff",
    86 => x"15555358",
    87 => x"a08082bc",
    88 => x"047b841d",
    89 => x"71087f5c",
    90 => x"555d5287",
    91 => x"56729c2a",
    92 => x"73842b54",
    93 => x"5271802e",
    94 => x"83388159",
    95 => x"b7125471",
    96 => x"89248438",
    97 => x"b0125478",
    98 => x"9438ff16",
    99 => x"56758025",
   100 => x"dc38800b",
   101 => x"ff115452",
   102 => x"a08082bc",
   103 => x"047351a0",
   104 => x"8083bd2d",
   105 => x"ff165675",
   106 => x"8025c238",
   107 => x"a0808392",
   108 => x"0477a080",
   109 => x"94f40c02",
   110 => x"80c0050d",
   111 => x"0402f805",
   112 => x"0d7352c0",
   113 => x"0870882a",
   114 => x"70810651",
   115 => x"51517080",
   116 => x"2ef13871",
   117 => x"c00c71a0",
   118 => x"8094f40c",
   119 => x"0288050d",
   120 => x"0402e805",
   121 => x"0d775675",
   122 => x"70840557",
   123 => x"08538054",
   124 => x"72982a73",
   125 => x"882b5452",
   126 => x"71802ea2",
   127 => x"38c00870",
   128 => x"882a7081",
   129 => x"06515151",
   130 => x"70802ef1",
   131 => x"3871c00c",
   132 => x"81158115",
   133 => x"55558374",
   134 => x"25d63871",
   135 => x"ca3874a0",
   136 => x"8094f40c",
   137 => x"0298050d",
   138 => x"0402f405",
   139 => x"0d747652",
   140 => x"53807125",
   141 => x"90387052",
   142 => x"72708405",
   143 => x"5408ff13",
   144 => x"535171f4",
   145 => x"38028c05",
   146 => x"0d0402d4",
   147 => x"050d7c7e",
   148 => x"5c58810b",
   149 => x"a0808ef8",
   150 => x"585a8359",
   151 => x"7608780c",
   152 => x"77087708",
   153 => x"56547375",
   154 => x"2e923877",
   155 => x"08537452",
   156 => x"a0808f88",
   157 => x"51a08080",
   158 => x"ed2d805a",
   159 => x"7756807b",
   160 => x"2590387a",
   161 => x"55757084",
   162 => x"055708ff",
   163 => x"16565474",
   164 => x"f4387708",
   165 => x"77085656",
   166 => x"75752e92",
   167 => x"38770853",
   168 => x"7452a080",
   169 => x"8fc851a0",
   170 => x"8080ed2d",
   171 => x"805aff19",
   172 => x"84185859",
   173 => x"788025ff",
   174 => x"a33879a0",
   175 => x"8094f40c",
   176 => x"02ac050d",
   177 => x"0402e405",
   178 => x"0d787a55",
   179 => x"56815785",
   180 => x"aad5aad5",
   181 => x"760cfad5",
   182 => x"aad5aa0b",
   183 => x"8c170ccc",
   184 => x"76a08080",
   185 => x"b92db30b",
   186 => x"8f17a080",
   187 => x"80b92d75",
   188 => x"085372fc",
   189 => x"e2d5aad5",
   190 => x"2e903875",
   191 => x"0852a080",
   192 => x"908851a0",
   193 => x"8080ed2d",
   194 => x"80578c16",
   195 => x"085574fa",
   196 => x"d5aad4b3",
   197 => x"2e91388c",
   198 => x"160852a0",
   199 => x"8090c451",
   200 => x"a08080ed",
   201 => x"2d805775",
   202 => x"55807425",
   203 => x"8e387470",
   204 => x"84055608",
   205 => x"ff155553",
   206 => x"73f43875",
   207 => x"085473fc",
   208 => x"e2d5aad5",
   209 => x"2e903875",
   210 => x"0852a080",
   211 => x"918051a0",
   212 => x"8080ed2d",
   213 => x"80578c16",
   214 => x"085372fa",
   215 => x"d5aad4b3",
   216 => x"2e91388c",
   217 => x"160852a0",
   218 => x"8091bc51",
   219 => x"a08080ed",
   220 => x"2d805776",
   221 => x"a08094f4",
   222 => x"0c029c05",
   223 => x"0d0402c4",
   224 => x"050d605b",
   225 => x"80629080",
   226 => x"8029ff05",
   227 => x"a08091f8",
   228 => x"53405aa0",
   229 => x"8080ed2d",
   230 => x"80e1b357",
   231 => x"80fe5eae",
   232 => x"51a08083",
   233 => x"bd2d7610",
   234 => x"70962a81",
   235 => x"06565774",
   236 => x"802e8538",
   237 => x"76810757",
   238 => x"76952a81",
   239 => x"06587780",
   240 => x"2e853876",
   241 => x"81325778",
   242 => x"77077f06",
   243 => x"775e598f",
   244 => x"ffff5876",
   245 => x"bfffff06",
   246 => x"707a3282",
   247 => x"2b7c1151",
   248 => x"57760c76",
   249 => x"1070962a",
   250 => x"81065657",
   251 => x"74802e85",
   252 => x"38768107",
   253 => x"5776952a",
   254 => x"81065574",
   255 => x"802e8538",
   256 => x"76813257",
   257 => x"ff185877",
   258 => x"8025c838",
   259 => x"7c578fff",
   260 => x"ff5876bf",
   261 => x"ffff0670",
   262 => x"7a32822b",
   263 => x"7c057008",
   264 => x"575e5674",
   265 => x"762e80e4",
   266 => x"38807a53",
   267 => x"a0809288",
   268 => x"525ca080",
   269 => x"80ed2d74",
   270 => x"54755375",
   271 => x"52a08092",
   272 => x"9c51a080",
   273 => x"80ed2d7b",
   274 => x"5a761070",
   275 => x"962a8106",
   276 => x"57577580",
   277 => x"2e853876",
   278 => x"81075776",
   279 => x"952a8106",
   280 => x"5574802e",
   281 => x"85387681",
   282 => x"3257ff18",
   283 => x"58778025",
   284 => x"ffa038ff",
   285 => x"1e5e7dfe",
   286 => x"a6388a51",
   287 => x"a08083bd",
   288 => x"2d7ba080",
   289 => x"94f40c02",
   290 => x"bc050d04",
   291 => x"811a5aa0",
   292 => x"8088c904",
   293 => x"02cc050d",
   294 => x"7e605e58",
   295 => x"815a805b",
   296 => x"80c07a58",
   297 => x"5c85ada9",
   298 => x"89bb780c",
   299 => x"79598156",
   300 => x"97557676",
   301 => x"07822b78",
   302 => x"11515485",
   303 => x"ada989bb",
   304 => x"740c7510",
   305 => x"ff165656",
   306 => x"748025e6",
   307 => x"38761081",
   308 => x"1a5a5798",
   309 => x"7925d738",
   310 => x"7756807d",
   311 => x"2590387c",
   312 => x"55757084",
   313 => x"055708ff",
   314 => x"16565474",
   315 => x"f4388157",
   316 => x"ff8787a5",
   317 => x"c3780c97",
   318 => x"5976822b",
   319 => x"78117008",
   320 => x"5f56567c",
   321 => x"ff8787a5",
   322 => x"c32e80c7",
   323 => x"38740854",
   324 => x"7385ada9",
   325 => x"89bb2e92",
   326 => x"38807508",
   327 => x"547653a0",
   328 => x"8092c452",
   329 => x"5aa08080",
   330 => x"ed2d7610",
   331 => x"ff1a5a57",
   332 => x"788025c5",
   333 => x"387a822b",
   334 => x"5675ad38",
   335 => x"7b52a080",
   336 => x"92e451a0",
   337 => x"8080ed2d",
   338 => x"7ba08094",
   339 => x"f40c02b4",
   340 => x"050d047a",
   341 => x"77077710",
   342 => x"ff1b5b58",
   343 => x"5b788025",
   344 => x"ff9738a0",
   345 => x"808ab504",
   346 => x"7552a080",
   347 => x"93a051a0",
   348 => x"8080ed2d",
   349 => x"75992a81",
   350 => x"32810670",
   351 => x"09810571",
   352 => x"07700970",
   353 => x"9f2c7d06",
   354 => x"79109fff",
   355 => x"fffc0660",
   356 => x"812a415a",
   357 => x"5d575859",
   358 => x"75da3879",
   359 => x"09810570",
   360 => x"7b079f2a",
   361 => x"55567bbf",
   362 => x"26843873",
   363 => x"9a388170",
   364 => x"53a08092",
   365 => x"e4525ca0",
   366 => x"8080ed2d",
   367 => x"7ba08094",
   368 => x"f40c02b4",
   369 => x"050d04a0",
   370 => x"8093b851",
   371 => x"a08080ed",
   372 => x"2d7b52a0",
   373 => x"8092e451",
   374 => x"a08080ed",
   375 => x"2d7ba080",
   376 => x"94f40c02",
   377 => x"b4050d04",
   378 => x"02dc050d",
   379 => x"810ba080",
   380 => x"8ef85858",
   381 => x"83597608",
   382 => x"800c8008",
   383 => x"77085654",
   384 => x"73752e92",
   385 => x"38800853",
   386 => x"7452a080",
   387 => x"8f8851a0",
   388 => x"8080ed2d",
   389 => x"80588070",
   390 => x"57557570",
   391 => x"84055708",
   392 => x"81165654",
   393 => x"a0807524",
   394 => x"f1388008",
   395 => x"77085656",
   396 => x"75752e92",
   397 => x"38800853",
   398 => x"7452a080",
   399 => x"8fc851a0",
   400 => x"8080ed2d",
   401 => x"8058ff19",
   402 => x"84185859",
   403 => x"788025ff",
   404 => x"a5387780",
   405 => x"2e8b38a0",
   406 => x"80948451",
   407 => x"a08080ed",
   408 => x"2d815785",
   409 => x"aad5aad5",
   410 => x"0b800cfa",
   411 => x"d5aad5aa",
   412 => x"0b8c0ccc",
   413 => x"0b800ba0",
   414 => x"8080b92d",
   415 => x"b30b8f0b",
   416 => x"a08080b9",
   417 => x"2d800855",
   418 => x"74fce2d5",
   419 => x"aad52e90",
   420 => x"38800852",
   421 => x"a0809088",
   422 => x"51a08080",
   423 => x"ed2d8057",
   424 => x"8c085877",
   425 => x"fad5aad4",
   426 => x"b32e9038",
   427 => x"8c0852a0",
   428 => x"8090c451",
   429 => x"a08080ed",
   430 => x"2d805780",
   431 => x"70575575",
   432 => x"70840557",
   433 => x"08811656",
   434 => x"54a08075",
   435 => x"24f13880",
   436 => x"085978fc",
   437 => x"e2d5aad5",
   438 => x"2e903880",
   439 => x"0852a080",
   440 => x"918051a0",
   441 => x"8080ed2d",
   442 => x"80578c08",
   443 => x"5473fad5",
   444 => x"aad4b32e",
   445 => x"80dd388c",
   446 => x"0852a080",
   447 => x"91bc51a0",
   448 => x"8080ed2d",
   449 => x"a0805280",
   450 => x"51a08089",
   451 => x"942da080",
   452 => x"94f40854",
   453 => x"a08094f4",
   454 => x"08802e8b",
   455 => x"38a08094",
   456 => x"a851a080",
   457 => x"80ed2d73",
   458 => x"528051a0",
   459 => x"8086fe2d",
   460 => x"a08094f4",
   461 => x"08802efd",
   462 => x"b338a080",
   463 => x"94c051a0",
   464 => x"8080ed2d",
   465 => x"810ba080",
   466 => x"8ef85858",
   467 => x"8359a080",
   468 => x"8bf60476",
   469 => x"802effac",
   470 => x"38a08094",
   471 => x"d851a080",
   472 => x"80ed2da0",
   473 => x"808e8404",
   474 => x"00ffffff",
   475 => x"ff00ffff",
   476 => x"ffff00ff",
   477 => x"ffffff00",
   478 => x"00000000",
   479 => x"55555555",
   480 => x"aaaaaaaa",
   481 => x"ffffffff",
   482 => x"53616e69",
   483 => x"74792063",
   484 => x"6865636b",
   485 => x"20666169",
   486 => x"6c656420",
   487 => x"28626566",
   488 => x"6f726520",
   489 => x"63616368",
   490 => x"65207265",
   491 => x"66726573",
   492 => x"6829206f",
   493 => x"6e203078",
   494 => x"25642028",
   495 => x"676f7420",
   496 => x"30782564",
   497 => x"290a0000",
   498 => x"53616e69",
   499 => x"74792063",
   500 => x"6865636b",
   501 => x"20666169",
   502 => x"6c656420",
   503 => x"28616674",
   504 => x"65722063",
   505 => x"61636865",
   506 => x"20726566",
   507 => x"72657368",
   508 => x"29206f6e",
   509 => x"20307825",
   510 => x"64202867",
   511 => x"6f742030",
   512 => x"78256429",
   513 => x"0a000000",
   514 => x"42797465",
   515 => x"20636865",
   516 => x"636b2066",
   517 => x"61696c65",
   518 => x"64202862",
   519 => x"65666f72",
   520 => x"65206361",
   521 => x"63686520",
   522 => x"72656672",
   523 => x"65736829",
   524 => x"20617420",
   525 => x"30202867",
   526 => x"6f742030",
   527 => x"78256429",
   528 => x"0a000000",
   529 => x"42797465",
   530 => x"20636865",
   531 => x"636b2066",
   532 => x"61696c65",
   533 => x"64202862",
   534 => x"65666f72",
   535 => x"65206361",
   536 => x"63686520",
   537 => x"72656672",
   538 => x"65736829",
   539 => x"20617420",
   540 => x"33202867",
   541 => x"6f742030",
   542 => x"78256429",
   543 => x"0a000000",
   544 => x"42797465",
   545 => x"20636865",
   546 => x"636b2066",
   547 => x"61696c65",
   548 => x"64202861",
   549 => x"66746572",
   550 => x"20636163",
   551 => x"68652072",
   552 => x"65667265",
   553 => x"73682920",
   554 => x"61742030",
   555 => x"2028676f",
   556 => x"74203078",
   557 => x"2564290a",
   558 => x"00000000",
   559 => x"42797465",
   560 => x"20636865",
   561 => x"636b2066",
   562 => x"61696c65",
   563 => x"64202861",
   564 => x"66746572",
   565 => x"20636163",
   566 => x"68652072",
   567 => x"65667265",
   568 => x"73682920",
   569 => x"61742033",
   570 => x"2028676f",
   571 => x"74203078",
   572 => x"2564290a",
   573 => x"00000000",
   574 => x"43686563",
   575 => x"6b696e67",
   576 => x"206d656d",
   577 => x"6f727900",
   578 => x"30782564",
   579 => x"20676f6f",
   580 => x"64207265",
   581 => x"6164732c",
   582 => x"20000000",
   583 => x"4572726f",
   584 => x"72206174",
   585 => x"20307825",
   586 => x"642c2065",
   587 => x"78706563",
   588 => x"74656420",
   589 => x"30782564",
   590 => x"2c20676f",
   591 => x"74203078",
   592 => x"25640a00",
   593 => x"42616420",
   594 => x"64617461",
   595 => x"20666f75",
   596 => x"6e642061",
   597 => x"74203078",
   598 => x"25642028",
   599 => x"30782564",
   600 => x"290a0000",
   601 => x"53445241",
   602 => x"4d207369",
   603 => x"7a652028",
   604 => x"61737375",
   605 => x"6d696e67",
   606 => x"206e6f20",
   607 => x"61646472",
   608 => x"65737320",
   609 => x"6661756c",
   610 => x"74732920",
   611 => x"69732030",
   612 => x"78256420",
   613 => x"6d656761",
   614 => x"62797465",
   615 => x"730a0000",
   616 => x"416c6961",
   617 => x"73657320",
   618 => x"666f756e",
   619 => x"64206174",
   620 => x"20307825",
   621 => x"640a0000",
   622 => x"28416c69",
   623 => x"61736573",
   624 => x"2070726f",
   625 => x"6261626c",
   626 => x"79207369",
   627 => x"6d706c79",
   628 => x"20696e64",
   629 => x"69636174",
   630 => x"65207468",
   631 => x"61742052",
   632 => x"414d0a69",
   633 => x"7320736d",
   634 => x"616c6c65",
   635 => x"72207468",
   636 => x"616e2036",
   637 => x"34206d65",
   638 => x"67616279",
   639 => x"74657329",
   640 => x"0a000000",
   641 => x"46697273",
   642 => x"74207374",
   643 => x"61676520",
   644 => x"73616e69",
   645 => x"74792063",
   646 => x"6865636b",
   647 => x"20706173",
   648 => x"7365642e",
   649 => x"0a000000",
   650 => x"41646472",
   651 => x"65737320",
   652 => x"63686563",
   653 => x"6b207061",
   654 => x"73736564",
   655 => x"2e0a0000",
   656 => x"4c465352",
   657 => x"20636865",
   658 => x"636b2070",
   659 => x"61737365",
   660 => x"642e0a0a",
   661 => x"00000000",
   662 => x"42797465",
   663 => x"20286471",
   664 => x"6d292063",
   665 => x"6865636b",
   666 => x"20706173",
   667 => x"7365640a",
   668 => x"00000000",
	others => x"00000000"
);

begin

process (clk)
begin
	if (clk'event and clk = '1') then
		if (from_zpu.memAWriteEnable = '1') and (from_zpu.memBWriteEnable = '1') and (from_zpu.memAAddr=from_zpu.memBAddr) and (from_zpu.memAWrite/=from_zpu.memBWrite) then
			report "write collision" severity failure;
		end if;
	
		if (from_zpu.memAWriteEnable = '1') then
			ram(to_integer(unsigned(from_zpu.memAAddr(maxAddrBit downto 2)))) := from_zpu.memAWrite;
			to_zpu.memARead <= from_zpu.memAWrite;
		else
			to_zpu.memARead <= ram(to_integer(unsigned(from_zpu.memAAddr(maxAddrBit downto 2))));
		end if;
	end if;
end process;

process (clk)
begin
	if (clk'event and clk = '1') then
		if (from_zpu.memBWriteEnable = '1') then
			ram(to_integer(unsigned(from_zpu.memBAddr(maxAddrBit downto 2)))) := from_zpu.memBWrite;
			to_zpu.memBRead <= from_zpu.memBWrite;
		else
			to_zpu.memBRead <= ram(to_integer(unsigned(from_zpu.memBAddr(maxAddrBit downto 2))));
		end if;
	end if;
end process;


end arch;

