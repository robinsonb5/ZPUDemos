-- ZPU
--
-- Copyright 2004-2008 oharboe - �yvind Harboe - oyvind.harboe@zylin.com
-- Modified by Alastair M. Robinson for the ZPUFlex project.
--
-- The FreeBSD license
-- 
-- Redistribution and use in source and binary forms, with or without
-- modification, are permitted provided that the following conditions
-- are met:
-- 
-- 1. Redistributions of source code must retain the above copyright
--    notice, this list of conditions and the following disclaimer.
-- 2. Redistributions in binary form must reproduce the above
--    copyright notice, this list of conditions and the following
--    disclaimer in the documentation and/or other materials
--    provided with the distribution.
-- 
-- THIS SOFTWARE IS PROVIDED BY THE ZPU PROJECT ``AS IS'' AND ANY
-- EXPRESS OR IMPLIED WARRANTIES, INCLUDING, BUT NOT LIMITED TO,
-- THE IMPLIED WARRANTIES OF MERCHANTABILITY AND FITNESS FOR A
-- PARTICULAR PURPOSE ARE DISCLAIMED. IN NO EVENT SHALL THE
-- ZPU PROJECT OR CONTRIBUTORS BE LIABLE FOR ANY DIRECT,
-- INDIRECT, INCIDENTAL, SPECIAL, EXEMPLARY, OR CONSEQUENTIAL DAMAGES
-- (INCLUDING, BUT NOT LIMITED TO, PROCUREMENT OF SUBSTITUTE GOODS
-- OR SERVICES; LOSS OF USE, DATA, OR PROFITS; OR BUSINESS INTERRUPTION)
-- HOWEVER CAUSED AND ON ANY THEORY OF LIABILITY, WHETHER IN CONTRACT,
-- STRICT LIABILITY, OR TORT (INCLUDING NEGLIGENCE OR OTHERWISE)
-- ARISING IN ANY WAY OUT OF THE USE OF THIS SOFTWARE, EVEN IF
-- ADVISED OF THE POSSIBILITY OF SUCH DAMAGE.
-- 
-- The views and conclusions contained in the software and documentation
-- are those of the authors and should not be interpreted as representing
-- official policies, either expressed or implied, of the ZPU Project.

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;


library work;
use work.zpu_config.all;
use work.zpupkg.all;

entity SDBootstrap_ROM is
generic
	(
		maxAddrBitBRAM : integer := maxAddrBitBRAMLimit -- Specify your actual ROM size to save LEs and unnecessary block RAM usage.
	);
port (
	clk : in std_logic;
	areset : in std_logic := '0';
	from_zpu : in ZPU_ToROM;
	to_zpu : out ZPU_FromROM
);
end SDBootstrap_ROM;

architecture arch of SDBootstrap_ROM is

type ram_type is array(natural range 0 to ((2**(maxAddrBitBRAM+1))/4)-1) of std_logic_vector(wordSize-1 downto 0);

shared variable ram : ram_type :=
(
     0 => x"84808080",
     1 => x"ee040000",
     2 => x"00000000",
     3 => x"84808080",
     4 => x"88080d80",
     5 => x"04848080",
     6 => x"80950471",
     7 => x"fd060872",
     8 => x"83060981",
     9 => x"05820583",
    10 => x"2b2a83ff",
    11 => x"ff065204",
    12 => x"71fc0608",
    13 => x"72830609",
    14 => x"81058305",
    15 => x"1010102a",
    16 => x"81ff0652",
    17 => x"0471fc06",
    18 => x"08848080",
    19 => x"a18c7383",
    20 => x"06101005",
    21 => x"08067381",
    22 => x"ff067383",
    23 => x"06098105",
    24 => x"83051010",
    25 => x"102b0772",
    26 => x"fc060c51",
    27 => x"51040284",
    28 => x"05848080",
    29 => x"80880c84",
    30 => x"80808095",
    31 => x"0b848080",
    32 => x"8e830400",
    33 => x"02c4050d",
    34 => x"0280c005",
    35 => x"83ffe0e0",
    36 => x"5b568076",
    37 => x"70840558",
    38 => x"08715e5e",
    39 => x"577c7084",
    40 => x"055e0858",
    41 => x"805b7798",
    42 => x"2a78882b",
    43 => x"59547389",
    44 => x"38765e84",
    45 => x"808083e3",
    46 => x"047b802e",
    47 => x"81fd3880",
    48 => x"5c7380e4",
    49 => x"2ea13873",
    50 => x"80e4268e",
    51 => x"387380e3",
    52 => x"2e819a38",
    53 => x"84808082",
    54 => x"fb047380",
    55 => x"f32e80f5",
    56 => x"38848080",
    57 => x"82fb0475",
    58 => x"84177108",
    59 => x"7e5c5557",
    60 => x"52728025",
    61 => x"8e38ad51",
    62 => x"84808083",
    63 => x"ee2d7209",
    64 => x"81055372",
    65 => x"802ebe38",
    66 => x"8755729c",
    67 => x"2a73842b",
    68 => x"54527180",
    69 => x"2e833881",
    70 => x"59897225",
    71 => x"8a38b712",
    72 => x"52848080",
    73 => x"82aa04b0",
    74 => x"12527880",
    75 => x"2e893871",
    76 => x"51848080",
    77 => x"83ee2dff",
    78 => x"15557480",
    79 => x"25cc3884",
    80 => x"808082cd",
    81 => x"04b05184",
    82 => x"808083ee",
    83 => x"2d805384",
    84 => x"80808394",
    85 => x"04758417",
    86 => x"71087054",
    87 => x"5c575284",
    88 => x"80808492",
    89 => x"2d7b5384",
    90 => x"80808394",
    91 => x"04758417",
    92 => x"71085657",
    93 => x"52848080",
    94 => x"83cb04a5",
    95 => x"51848080",
    96 => x"83ee2d73",
    97 => x"51848080",
    98 => x"83ee2d82",
    99 => x"17578480",
   100 => x"8083d604",
   101 => x"72ff1454",
   102 => x"52807225",
   103 => x"b9387970",
   104 => x"81055b84",
   105 => x"808080b0",
   106 => x"2d705254",
   107 => x"84808083",
   108 => x"ee2d8117",
   109 => x"57848080",
   110 => x"83940473",
   111 => x"a52e0981",
   112 => x"06893881",
   113 => x"5c848080",
   114 => x"83d60473",
   115 => x"51848080",
   116 => x"83ee2d81",
   117 => x"1757811b",
   118 => x"5b837b25",
   119 => x"fdc83873",
   120 => x"fdbb387d",
   121 => x"83ffe080",
   122 => x"0c02bc05",
   123 => x"0d0402f8",
   124 => x"050d7352",
   125 => x"c0087088",
   126 => x"2a708106",
   127 => x"51515170",
   128 => x"802ef138",
   129 => x"71c00c71",
   130 => x"83ffe080",
   131 => x"0c028805",
   132 => x"0d0402e8",
   133 => x"050d8078",
   134 => x"57557570",
   135 => x"84055708",
   136 => x"53805472",
   137 => x"982a7388",
   138 => x"2b545271",
   139 => x"802ea238",
   140 => x"c0087088",
   141 => x"2a708106",
   142 => x"51515170",
   143 => x"802ef138",
   144 => x"71c00c81",
   145 => x"15811555",
   146 => x"55837425",
   147 => x"d63871ca",
   148 => x"387483ff",
   149 => x"e0800c02",
   150 => x"98050d04",
   151 => x"02f4050d",
   152 => x"d45281ff",
   153 => x"720c7108",
   154 => x"5381ff72",
   155 => x"0c72882b",
   156 => x"83fe8006",
   157 => x"72087081",
   158 => x"ff065152",
   159 => x"5381ff72",
   160 => x"0c727107",
   161 => x"882b7208",
   162 => x"7081ff06",
   163 => x"51525381",
   164 => x"ff720c72",
   165 => x"7107882b",
   166 => x"72087081",
   167 => x"ff067207",
   168 => x"83ffe080",
   169 => x"0c525302",
   170 => x"8c050d04",
   171 => x"02f4050d",
   172 => x"74767181",
   173 => x"ff06d40c",
   174 => x"535383ff",
   175 => x"f1a00885",
   176 => x"3871892b",
   177 => x"5271982a",
   178 => x"d40c7190",
   179 => x"2a7081ff",
   180 => x"06d40c51",
   181 => x"71882a70",
   182 => x"81ff06d4",
   183 => x"0c517181",
   184 => x"ff06d40c",
   185 => x"72902a70",
   186 => x"81ff06d4",
   187 => x"0c51d408",
   188 => x"7081ff06",
   189 => x"515182b8",
   190 => x"bf527081",
   191 => x"ff2e0981",
   192 => x"06943881",
   193 => x"ff0bd40c",
   194 => x"d4087081",
   195 => x"ff06ff14",
   196 => x"54515171",
   197 => x"e5387083",
   198 => x"ffe0800c",
   199 => x"028c050d",
   200 => x"0402fc05",
   201 => x"0d81c751",
   202 => x"81ff0bd4",
   203 => x"0cff1151",
   204 => x"708025f4",
   205 => x"38028405",
   206 => x"0d0402f0",
   207 => x"050d8480",
   208 => x"8086a12d",
   209 => x"819c9f53",
   210 => x"805287fc",
   211 => x"80f75184",
   212 => x"808085ac",
   213 => x"2d83ffe0",
   214 => x"80085483",
   215 => x"ffe08008",
   216 => x"812e0981",
   217 => x"06ae3881",
   218 => x"ff0bd40c",
   219 => x"820a5284",
   220 => x"9c80e951",
   221 => x"84808085",
   222 => x"ac2d83ff",
   223 => x"e080088e",
   224 => x"3881ff0b",
   225 => x"d40c7353",
   226 => x"84808087",
   227 => x"9b048480",
   228 => x"8086a12d",
   229 => x"ff135372",
   230 => x"ffae3872",
   231 => x"83ffe080",
   232 => x"0c029005",
   233 => x"0d0402f4",
   234 => x"050d81ff",
   235 => x"0bd40c84",
   236 => x"8080a19c",
   237 => x"51848080",
   238 => x"84922d93",
   239 => x"53805287",
   240 => x"fc80c151",
   241 => x"84808085",
   242 => x"ac2d83ff",
   243 => x"e080088e",
   244 => x"3881ff0b",
   245 => x"d40c8153",
   246 => x"84808087",
   247 => x"ea048480",
   248 => x"8086a12d",
   249 => x"ff135372",
   250 => x"d4387283",
   251 => x"ffe0800c",
   252 => x"028c050d",
   253 => x"0402f005",
   254 => x"0d848080",
   255 => x"86a12d83",
   256 => x"aa52849c",
   257 => x"80c85184",
   258 => x"808085ac",
   259 => x"2d83ffe0",
   260 => x"800883ff",
   261 => x"e0800853",
   262 => x"848080a1",
   263 => x"a8525384",
   264 => x"80808184",
   265 => x"2d72812e",
   266 => x"098106a9",
   267 => x"38848080",
   268 => x"84dc2d83",
   269 => x"ffe08008",
   270 => x"83ffff06",
   271 => x"537283aa",
   272 => x"2ebb3883",
   273 => x"ffe08008",
   274 => x"52848080",
   275 => x"a1c05184",
   276 => x"80808184",
   277 => x"2d848080",
   278 => x"87a62d84",
   279 => x"808088f5",
   280 => x"04815484",
   281 => x"80808aa0",
   282 => x"04848080",
   283 => x"a1d85184",
   284 => x"80808184",
   285 => x"2d805484",
   286 => x"80808aa0",
   287 => x"0481ff0b",
   288 => x"d40cb153",
   289 => x"84808086",
   290 => x"ba2d83ff",
   291 => x"e0800880",
   292 => x"2e80fe38",
   293 => x"805287fc",
   294 => x"80fa5184",
   295 => x"808085ac",
   296 => x"2d83ffe0",
   297 => x"800880d7",
   298 => x"3883ffe0",
   299 => x"80085284",
   300 => x"8080a1f4",
   301 => x"51848080",
   302 => x"81842d81",
   303 => x"ff0bd40c",
   304 => x"d4087081",
   305 => x"ff067054",
   306 => x"848080a2",
   307 => x"80535153",
   308 => x"84808081",
   309 => x"842d81ff",
   310 => x"0bd40c81",
   311 => x"ff0bd40c",
   312 => x"81ff0bd4",
   313 => x"0c81ff0b",
   314 => x"d40c7286",
   315 => x"2a708106",
   316 => x"70565153",
   317 => x"72802ea8",
   318 => x"38848080",
   319 => x"88e10483",
   320 => x"ffe08008",
   321 => x"52848080",
   322 => x"a1f45184",
   323 => x"80808184",
   324 => x"2d72822e",
   325 => x"fed338ff",
   326 => x"135372fe",
   327 => x"e7387254",
   328 => x"7383ffe0",
   329 => x"800c0290",
   330 => x"050d0402",
   331 => x"f4050d81",
   332 => x"0b83fff1",
   333 => x"a00cd008",
   334 => x"708f2a70",
   335 => x"81065151",
   336 => x"5372f338",
   337 => x"72d00c84",
   338 => x"808086a1",
   339 => x"2dd00870",
   340 => x"8f2a7081",
   341 => x"06515153",
   342 => x"72f33881",
   343 => x"0bd00c87",
   344 => x"53805284",
   345 => x"d480c051",
   346 => x"84808085",
   347 => x"ac2d83ff",
   348 => x"e0800881",
   349 => x"2e973872",
   350 => x"822e0981",
   351 => x"06893880",
   352 => x"53848080",
   353 => x"8bc704ff",
   354 => x"135372d5",
   355 => x"38848080",
   356 => x"87f52d83",
   357 => x"ffe08008",
   358 => x"83fff1a0",
   359 => x"0c815287",
   360 => x"fc80d051",
   361 => x"84808085",
   362 => x"ac2d81ff",
   363 => x"0bd40cd0",
   364 => x"08708f2a",
   365 => x"70810651",
   366 => x"515372f3",
   367 => x"3872d00c",
   368 => x"81ff0bd4",
   369 => x"0c815372",
   370 => x"83ffe080",
   371 => x"0c028c05",
   372 => x"0d04800b",
   373 => x"83ffe080",
   374 => x"0c0402e0",
   375 => x"050d797b",
   376 => x"57578058",
   377 => x"81ff0bd4",
   378 => x"0cd00870",
   379 => x"8f2a7081",
   380 => x"06515154",
   381 => x"73f33882",
   382 => x"810bd00c",
   383 => x"81ff0bd4",
   384 => x"0c765287",
   385 => x"fc80d151",
   386 => x"84808085",
   387 => x"ac2d80db",
   388 => x"c6df5583",
   389 => x"ffe08008",
   390 => x"802e9b38",
   391 => x"83ffe080",
   392 => x"08537652",
   393 => x"848080a2",
   394 => x"90518480",
   395 => x"8081842d",
   396 => x"8480808d",
   397 => x"8c0481ff",
   398 => x"0bd40cd4",
   399 => x"087081ff",
   400 => x"06515473",
   401 => x"81fe2e09",
   402 => x"8106a538",
   403 => x"80ff5484",
   404 => x"808084dc",
   405 => x"2d83ffe0",
   406 => x"80087670",
   407 => x"8405580c",
   408 => x"ff145473",
   409 => x"8025e838",
   410 => x"81588480",
   411 => x"808cf604",
   412 => x"ff155574",
   413 => x"c13881ff",
   414 => x"0bd40cd0",
   415 => x"08708f2a",
   416 => x"70810651",
   417 => x"515473f3",
   418 => x"3873d00c",
   419 => x"7783ffe0",
   420 => x"800c02a0",
   421 => x"050d0402",
   422 => x"f4050d74",
   423 => x"70882a83",
   424 => x"fe800670",
   425 => x"72982a07",
   426 => x"72882b87",
   427 => x"fc808006",
   428 => x"73982b81",
   429 => x"f00a0671",
   430 => x"73070783",
   431 => x"ffe0800c",
   432 => x"56515351",
   433 => x"028c050d",
   434 => x"0402f805",
   435 => x"0d028e05",
   436 => x"84808080",
   437 => x"b02d7498",
   438 => x"2b71902b",
   439 => x"0770902c",
   440 => x"83ffe080",
   441 => x"0c525202",
   442 => x"88050d04",
   443 => x"02f8050d",
   444 => x"7370902b",
   445 => x"71902a07",
   446 => x"83ffe080",
   447 => x"0c520288",
   448 => x"050d0402",
   449 => x"ec050d80",
   450 => x"0bfc800c",
   451 => x"848080a2",
   452 => x"b0518480",
   453 => x"8084922d",
   454 => x"8480808a",
   455 => x"ab2d83ff",
   456 => x"e0800880",
   457 => x"2e828638",
   458 => x"848080a2",
   459 => x"c8518480",
   460 => x"8084922d",
   461 => x"84808091",
   462 => x"912d83ff",
   463 => x"e1a05284",
   464 => x"8080a2e0",
   465 => x"51848080",
   466 => x"9df42d83",
   467 => x"ffe08008",
   468 => x"802e81cd",
   469 => x"3883ffe1",
   470 => x"a00b8480",
   471 => x"80a2ec52",
   472 => x"54848080",
   473 => x"84922d80",
   474 => x"55737081",
   475 => x"05558480",
   476 => x"8080b02d",
   477 => x"5372a02e",
   478 => x"80e63872",
   479 => x"c00c72a3",
   480 => x"2e818438",
   481 => x"7280c72e",
   482 => x"0981068d",
   483 => x"38848080",
   484 => x"808c2d84",
   485 => x"80808fbb",
   486 => x"04728a2e",
   487 => x"0981068d",
   488 => x"38848080",
   489 => x"80952d84",
   490 => x"80808fbb",
   491 => x"047280cc",
   492 => x"2e098106",
   493 => x"863883ff",
   494 => x"e1a05472",
   495 => x"81df06f0",
   496 => x"057081ff",
   497 => x"065153b8",
   498 => x"73278938",
   499 => x"ef137081",
   500 => x"ff065153",
   501 => x"74842b73",
   502 => x"07558480",
   503 => x"808ee904",
   504 => x"72a32ea3",
   505 => x"38737081",
   506 => x"05558480",
   507 => x"8080b02d",
   508 => x"5372a02e",
   509 => x"f038ff14",
   510 => x"75537052",
   511 => x"54848080",
   512 => x"9df42d74",
   513 => x"fc800c73",
   514 => x"70810555",
   515 => x"84808080",
   516 => x"b02d5372",
   517 => x"8a2e0981",
   518 => x"06ed3884",
   519 => x"80808ee7",
   520 => x"04848080",
   521 => x"a3805184",
   522 => x"80808492",
   523 => x"2d848080",
   524 => x"a39c5184",
   525 => x"80808492",
   526 => x"2d800b83",
   527 => x"ffe0800c",
   528 => x"0294050d",
   529 => x"0402e805",
   530 => x"0d77797b",
   531 => x"58555580",
   532 => x"53727625",
   533 => x"af387470",
   534 => x"81055684",
   535 => x"808080b0",
   536 => x"2d747081",
   537 => x"05568480",
   538 => x"8080b02d",
   539 => x"52527171",
   540 => x"2e893881",
   541 => x"51848080",
   542 => x"91860481",
   543 => x"13538480",
   544 => x"8090d104",
   545 => x"80517083",
   546 => x"ffe0800c",
   547 => x"0298050d",
   548 => x"0402d805",
   549 => x"0dff0b83",
   550 => x"fff5cc0c",
   551 => x"800b83ff",
   552 => x"f5e00c84",
   553 => x"8080a3a8",
   554 => x"51848080",
   555 => x"84922d83",
   556 => x"fff1b852",
   557 => x"80518480",
   558 => x"808bda2d",
   559 => x"83ffe080",
   560 => x"085483ff",
   561 => x"e0800895",
   562 => x"38848080",
   563 => x"a3b85184",
   564 => x"80808492",
   565 => x"2d735584",
   566 => x"808099b6",
   567 => x"04848080",
   568 => x"a3cc5184",
   569 => x"80808492",
   570 => x"2d805681",
   571 => x"0b83fff1",
   572 => x"ac0c8853",
   573 => x"848080a3",
   574 => x"e45283ff",
   575 => x"f1ee5184",
   576 => x"808090c5",
   577 => x"2d83ffe0",
   578 => x"8008762e",
   579 => x"0981068b",
   580 => x"3883ffe0",
   581 => x"800883ff",
   582 => x"f1ac0c88",
   583 => x"53848080",
   584 => x"a3f05283",
   585 => x"fff28a51",
   586 => x"84808090",
   587 => x"c52d83ff",
   588 => x"e080088b",
   589 => x"3883ffe0",
   590 => x"800883ff",
   591 => x"f1ac0c83",
   592 => x"fff1ac08",
   593 => x"52848080",
   594 => x"a3fc5184",
   595 => x"80808184",
   596 => x"2d83fff1",
   597 => x"ac08802e",
   598 => x"81cb3883",
   599 => x"fff4fe0b",
   600 => x"84808080",
   601 => x"b02d83ff",
   602 => x"f4ff0b84",
   603 => x"808080b0",
   604 => x"2d71982b",
   605 => x"71902b07",
   606 => x"83fff580",
   607 => x"0b848080",
   608 => x"80b02d70",
   609 => x"882b7207",
   610 => x"83fff581",
   611 => x"0b848080",
   612 => x"80b02d71",
   613 => x"0783fff5",
   614 => x"b60b8480",
   615 => x"8080b02d",
   616 => x"83fff5b7",
   617 => x"0b848080",
   618 => x"80b02d71",
   619 => x"882b0753",
   620 => x"5f54525a",
   621 => x"56575573",
   622 => x"81abaa2e",
   623 => x"09810695",
   624 => x"38755184",
   625 => x"80808d97",
   626 => x"2d83ffe0",
   627 => x"80085684",
   628 => x"808093ee",
   629 => x"047382d4",
   630 => x"d52e9338",
   631 => x"848080a4",
   632 => x"90518480",
   633 => x"8084922d",
   634 => x"84808095",
   635 => x"fa047552",
   636 => x"848080a4",
   637 => x"b0518480",
   638 => x"8081842d",
   639 => x"83fff1b8",
   640 => x"52755184",
   641 => x"80808bda",
   642 => x"2d83ffe0",
   643 => x"80085583",
   644 => x"ffe08008",
   645 => x"802e859e",
   646 => x"38848080",
   647 => x"a4c85184",
   648 => x"80808492",
   649 => x"2d848080",
   650 => x"a4f05184",
   651 => x"80808184",
   652 => x"2d885384",
   653 => x"8080a3f0",
   654 => x"5283fff2",
   655 => x"8a518480",
   656 => x"8090c52d",
   657 => x"83ffe080",
   658 => x"088e3881",
   659 => x"0b83fff5",
   660 => x"e00c8480",
   661 => x"80958604",
   662 => x"88538480",
   663 => x"80a3e452",
   664 => x"83fff1ee",
   665 => x"51848080",
   666 => x"90c52d83",
   667 => x"ffe08008",
   668 => x"802e9338",
   669 => x"848080a5",
   670 => x"88518480",
   671 => x"8081842d",
   672 => x"84808095",
   673 => x"fa0483ff",
   674 => x"f5b60b84",
   675 => x"808080b0",
   676 => x"2d547380",
   677 => x"d52e0981",
   678 => x"0680df38",
   679 => x"83fff5b7",
   680 => x"0b848080",
   681 => x"80b02d54",
   682 => x"7381aa2e",
   683 => x"09810680",
   684 => x"c938800b",
   685 => x"83fff1b8",
   686 => x"0b848080",
   687 => x"80b02d56",
   688 => x"547481e9",
   689 => x"2e833881",
   690 => x"547481eb",
   691 => x"2e8c3880",
   692 => x"5573752e",
   693 => x"09810683",
   694 => x"dd3883ff",
   695 => x"f1c30b84",
   696 => x"808080b0",
   697 => x"2d557492",
   698 => x"3883fff1",
   699 => x"c40b8480",
   700 => x"8080b02d",
   701 => x"5473822e",
   702 => x"89388055",
   703 => x"84808099",
   704 => x"b60483ff",
   705 => x"f1c50b84",
   706 => x"808080b0",
   707 => x"2d7083ff",
   708 => x"f5e80cff",
   709 => x"0583fff5",
   710 => x"dc0c83ff",
   711 => x"f1c60b84",
   712 => x"808080b0",
   713 => x"2d83fff1",
   714 => x"c70b8480",
   715 => x"8080b02d",
   716 => x"58760577",
   717 => x"82802905",
   718 => x"7083fff5",
   719 => x"d00c83ff",
   720 => x"f1c80b84",
   721 => x"808080b0",
   722 => x"2d7083ff",
   723 => x"f5c80c83",
   724 => x"fff5e008",
   725 => x"59575876",
   726 => x"802e81ea",
   727 => x"38885384",
   728 => x"8080a3f0",
   729 => x"5283fff2",
   730 => x"8a518480",
   731 => x"8090c52d",
   732 => x"83ffe080",
   733 => x"0882bf38",
   734 => x"83fff5e8",
   735 => x"0870842b",
   736 => x"83fff5b8",
   737 => x"0c7083ff",
   738 => x"f5e40c83",
   739 => x"fff1dd0b",
   740 => x"84808080",
   741 => x"b02d83ff",
   742 => x"f1dc0b84",
   743 => x"808080b0",
   744 => x"2d718280",
   745 => x"290583ff",
   746 => x"f1de0b84",
   747 => x"808080b0",
   748 => x"2d708480",
   749 => x"80291283",
   750 => x"fff1df0b",
   751 => x"84808080",
   752 => x"b02d7081",
   753 => x"800a2912",
   754 => x"7083fff1",
   755 => x"b00c83ff",
   756 => x"f5c80871",
   757 => x"2983fff5",
   758 => x"d0080570",
   759 => x"83fff5f0",
   760 => x"0c83fff1",
   761 => x"e50b8480",
   762 => x"8080b02d",
   763 => x"83fff1e4",
   764 => x"0b848080",
   765 => x"80b02d71",
   766 => x"82802905",
   767 => x"83fff1e6",
   768 => x"0b848080",
   769 => x"80b02d70",
   770 => x"84808029",
   771 => x"1283fff1",
   772 => x"e70b8480",
   773 => x"8080b02d",
   774 => x"70982b81",
   775 => x"f00a0672",
   776 => x"057083ff",
   777 => x"f1b40cfe",
   778 => x"117e2977",
   779 => x"0583fff5",
   780 => x"d80c5259",
   781 => x"5243545e",
   782 => x"51525952",
   783 => x"5d575957",
   784 => x"84808099",
   785 => x"b40483ff",
   786 => x"f1ca0b84",
   787 => x"808080b0",
   788 => x"2d83fff1",
   789 => x"c90b8480",
   790 => x"8080b02d",
   791 => x"71828029",
   792 => x"057083ff",
   793 => x"f5b80c70",
   794 => x"a02983ff",
   795 => x"0570892a",
   796 => x"7083fff5",
   797 => x"e40c83ff",
   798 => x"f1cf0b84",
   799 => x"808080b0",
   800 => x"2d83fff1",
   801 => x"ce0b8480",
   802 => x"8080b02d",
   803 => x"71828029",
   804 => x"057083ff",
   805 => x"f1b00c7b",
   806 => x"71291e70",
   807 => x"83fff5d8",
   808 => x"0c7d83ff",
   809 => x"f1b40c73",
   810 => x"0583fff5",
   811 => x"f00c555e",
   812 => x"51515555",
   813 => x"81557483",
   814 => x"ffe0800c",
   815 => x"02a8050d",
   816 => x"0402ec05",
   817 => x"0d767087",
   818 => x"2c7180ff",
   819 => x"06575553",
   820 => x"83fff5e0",
   821 => x"088a3872",
   822 => x"882c7381",
   823 => x"ff065654",
   824 => x"7383fff5",
   825 => x"cc082ea9",
   826 => x"3883fff1",
   827 => x"b85283ff",
   828 => x"f5d00814",
   829 => x"51848080",
   830 => x"8bda2d83",
   831 => x"ffe08008",
   832 => x"5383ffe0",
   833 => x"8008802e",
   834 => x"80cf3873",
   835 => x"83fff5cc",
   836 => x"0c83fff5",
   837 => x"e008802e",
   838 => x"a2387484",
   839 => x"2983fff1",
   840 => x"b8057008",
   841 => x"52538480",
   842 => x"808d972d",
   843 => x"83ffe080",
   844 => x"08f00a06",
   845 => x"55848080",
   846 => x"9ad70474",
   847 => x"1083fff1",
   848 => x"b8057084",
   849 => x"8080809b",
   850 => x"2d525384",
   851 => x"80808dc9",
   852 => x"2d83ffe0",
   853 => x"80085574",
   854 => x"537283ff",
   855 => x"e0800c02",
   856 => x"94050d04",
   857 => x"02cc050d",
   858 => x"7e605e5b",
   859 => x"8056ff0b",
   860 => x"83fff5cc",
   861 => x"0c83fff1",
   862 => x"b40883ff",
   863 => x"f5d80856",
   864 => x"5783fff5",
   865 => x"e008762e",
   866 => x"8f3883ff",
   867 => x"f5e80884",
   868 => x"2b598480",
   869 => x"809ba004",
   870 => x"83fff5e4",
   871 => x"08842b59",
   872 => x"805a7979",
   873 => x"2781f038",
   874 => x"798f06a0",
   875 => x"17575473",
   876 => x"a4387452",
   877 => x"848080a5",
   878 => x"a8518480",
   879 => x"8081842d",
   880 => x"83fff1b8",
   881 => x"52745181",
   882 => x"15558480",
   883 => x"808bda2d",
   884 => x"83fff1b8",
   885 => x"56807684",
   886 => x"808080b0",
   887 => x"2d555873",
   888 => x"782e8338",
   889 => x"81587381",
   890 => x"e52e81a2",
   891 => x"38817079",
   892 => x"06555c73",
   893 => x"802e8196",
   894 => x"388b1684",
   895 => x"808080b0",
   896 => x"2d980658",
   897 => x"77818738",
   898 => x"8b537c52",
   899 => x"75518480",
   900 => x"8090c52d",
   901 => x"83ffe080",
   902 => x"0880f338",
   903 => x"9c160851",
   904 => x"8480808d",
   905 => x"972d83ff",
   906 => x"e0800884",
   907 => x"1c0c9a16",
   908 => x"84808080",
   909 => x"9b2d5184",
   910 => x"80808dc9",
   911 => x"2d83ffe0",
   912 => x"800883ff",
   913 => x"e0800855",
   914 => x"5583fff5",
   915 => x"e008802e",
   916 => x"a0389416",
   917 => x"84808080",
   918 => x"9b2d5184",
   919 => x"80808dc9",
   920 => x"2d83ffe0",
   921 => x"8008902b",
   922 => x"83fff00a",
   923 => x"06701651",
   924 => x"5473881c",
   925 => x"0c777b0c",
   926 => x"7c528480",
   927 => x"80a5c851",
   928 => x"84808081",
   929 => x"842d7b54",
   930 => x"8480809d",
   931 => x"e904811a",
   932 => x"5a848080",
   933 => x"9ba20483",
   934 => x"fff5e008",
   935 => x"802e80c7",
   936 => x"38765184",
   937 => x"808099c1",
   938 => x"2d83ffe0",
   939 => x"800883ff",
   940 => x"e0800853",
   941 => x"848080a5",
   942 => x"dc525784",
   943 => x"80808184",
   944 => x"2d7680ff",
   945 => x"fffff806",
   946 => x"547380ff",
   947 => x"fffff82e",
   948 => x"9638fe17",
   949 => x"83fff5e8",
   950 => x"082983ff",
   951 => x"f5f00805",
   952 => x"55848080",
   953 => x"9ba00480",
   954 => x"547383ff",
   955 => x"e0800c02",
   956 => x"b4050d04",
   957 => x"02d4050d",
   958 => x"7c7e7154",
   959 => x"83fff5bc",
   960 => x"535a5784",
   961 => x"80809ae4",
   962 => x"2d83ffe0",
   963 => x"800881ff",
   964 => x"06567580",
   965 => x"2e81b938",
   966 => x"848080a5",
   967 => x"f4518480",
   968 => x"8084922d",
   969 => x"83fff5c0",
   970 => x"0883ff05",
   971 => x"892a5b80",
   972 => x"70595a79",
   973 => x"7b2581b8",
   974 => x"3883fff5",
   975 => x"c408fe11",
   976 => x"83fff5e8",
   977 => x"082983ff",
   978 => x"f5f00811",
   979 => x"7a83fff5",
   980 => x"dc080605",
   981 => x"7a585157",
   982 => x"5483fff5",
   983 => x"f0085375",
   984 => x"52848080",
   985 => x"a6905184",
   986 => x"80808184",
   987 => x"2d785275",
   988 => x"51848080",
   989 => x"8bda2d83",
   990 => x"ffe08008",
   991 => x"802e80e4",
   992 => x"38848080",
   993 => x"a6b45184",
   994 => x"80808492",
   995 => x"2d811870",
   996 => x"83fff5dc",
   997 => x"08065758",
   998 => x"75a33884",
   999 => x"8080a6c4",
  1000 => x"51848080",
  1001 => x"84922d83",
  1002 => x"fff5c408",
  1003 => x"51848080",
  1004 => x"99c12d83",
  1005 => x"ffe08008",
  1006 => x"83fff5c4",
  1007 => x"0c848019",
  1008 => x"811b5b59",
  1009 => x"7a7a24fe",
  1010 => x"f0388480",
  1011 => x"809ff004",
  1012 => x"76528480",
  1013 => x"80a6dc51",
  1014 => x"84808081",
  1015 => x"842d8480",
  1016 => x"809ff204",
  1017 => x"83ffe080",
  1018 => x"08568480",
  1019 => x"809ff204",
  1020 => x"81567583",
  1021 => x"ffe0800c",
  1022 => x"02ac050d",
  1023 => x"0483ffe0",
  1024 => x"8c080283",
  1025 => x"ffe08c0c",
  1026 => x"ff3d0d80",
  1027 => x"0b83ffe0",
  1028 => x"8c08fc05",
  1029 => x"0c83ffe0",
  1030 => x"8c088805",
  1031 => x"088106ff",
  1032 => x"11700970",
  1033 => x"83ffe08c",
  1034 => x"088c0508",
  1035 => x"0683ffe0",
  1036 => x"8c08fc05",
  1037 => x"081183ff",
  1038 => x"e08c08fc",
  1039 => x"050c83ff",
  1040 => x"e08c0888",
  1041 => x"0508812a",
  1042 => x"83ffe08c",
  1043 => x"0888050c",
  1044 => x"83ffe08c",
  1045 => x"088c0508",
  1046 => x"1083ffe0",
  1047 => x"8c088c05",
  1048 => x"0c515151",
  1049 => x"5183ffe0",
  1050 => x"8c088805",
  1051 => x"08802e84",
  1052 => x"38ffa239",
  1053 => x"83ffe08c",
  1054 => x"08fc0508",
  1055 => x"7083ffe0",
  1056 => x"800c5183",
  1057 => x"3d0d83ff",
  1058 => x"e08c0c04",
  1059 => x"00ffffff",
  1060 => x"ff00ffff",
  1061 => x"ffff00ff",
  1062 => x"ffffff00",
  1063 => x"436d645f",
  1064 => x"696e6974",
  1065 => x"0a000000",
  1066 => x"636d645f",
  1067 => x"434d4438",
  1068 => x"20726573",
  1069 => x"706f6e73",
  1070 => x"653a2025",
  1071 => x"640a0000",
  1072 => x"434d4438",
  1073 => x"5f342072",
  1074 => x"6573706f",
  1075 => x"6e73653a",
  1076 => x"2025640a",
  1077 => x"00000000",
  1078 => x"53444843",
  1079 => x"20496e69",
  1080 => x"7469616c",
  1081 => x"697a6174",
  1082 => x"696f6e20",
  1083 => x"6572726f",
  1084 => x"72210a00",
  1085 => x"434d4435",
  1086 => x"38202564",
  1087 => x"0a202000",
  1088 => x"434d4435",
  1089 => x"385f3220",
  1090 => x"25640a20",
  1091 => x"20000000",
  1092 => x"52656164",
  1093 => x"20636f6d",
  1094 => x"6d616e64",
  1095 => x"20666169",
  1096 => x"6c656420",
  1097 => x"61742025",
  1098 => x"64202825",
  1099 => x"64290a00",
  1100 => x"496e6974",
  1101 => x"69616c69",
  1102 => x"7a696e67",
  1103 => x"20534420",
  1104 => x"63617264",
  1105 => x"0a000000",
  1106 => x"48756e74",
  1107 => x"696e6720",
  1108 => x"666f7220",
  1109 => x"70617274",
  1110 => x"6974696f",
  1111 => x"6e0a0000",
  1112 => x"4d414e49",
  1113 => x"46455354",
  1114 => x"4d535400",
  1115 => x"50617273",
  1116 => x"696e6720",
  1117 => x"6d616e69",
  1118 => x"66657374",
  1119 => x"0a000000",
  1120 => x"4c6f6164",
  1121 => x"696e6720",
  1122 => x"6d616e69",
  1123 => x"66657374",
  1124 => x"20666169",
  1125 => x"6c65640a",
  1126 => x"00000000",
  1127 => x"52657475",
  1128 => x"726e696e",
  1129 => x"670a0000",
  1130 => x"52656164",
  1131 => x"696e6720",
  1132 => x"4d42520a",
  1133 => x"00000000",
  1134 => x"52656164",
  1135 => x"206f6620",
  1136 => x"4d425220",
  1137 => x"6661696c",
  1138 => x"65640a00",
  1139 => x"4d425220",
  1140 => x"73756363",
  1141 => x"65737366",
  1142 => x"756c6c79",
  1143 => x"20726561",
  1144 => x"640a0000",
  1145 => x"46415431",
  1146 => x"36202020",
  1147 => x"00000000",
  1148 => x"46415433",
  1149 => x"32202020",
  1150 => x"00000000",
  1151 => x"50617274",
  1152 => x"6974696f",
  1153 => x"6e636f75",
  1154 => x"6e742025",
  1155 => x"640a0000",
  1156 => x"4e6f2070",
  1157 => x"61727469",
  1158 => x"74696f6e",
  1159 => x"20736967",
  1160 => x"6e617475",
  1161 => x"72652066",
  1162 => x"6f756e64",
  1163 => x"0a000000",
  1164 => x"52656164",
  1165 => x"696e6720",
  1166 => x"626f6f74",
  1167 => x"20736563",
  1168 => x"746f7220",
  1169 => x"25640a00",
  1170 => x"52656164",
  1171 => x"20626f6f",
  1172 => x"74207365",
  1173 => x"63746f72",
  1174 => x"2066726f",
  1175 => x"6d206669",
  1176 => x"72737420",
  1177 => x"70617274",
  1178 => x"6974696f",
  1179 => x"6e0a0000",
  1180 => x"48756e74",
  1181 => x"696e6720",
  1182 => x"666f7220",
  1183 => x"66696c65",
  1184 => x"73797374",
  1185 => x"656d0a00",
  1186 => x"556e7375",
  1187 => x"70706f72",
  1188 => x"74656420",
  1189 => x"70617274",
  1190 => x"6974696f",
  1191 => x"6e207479",
  1192 => x"7065210d",
  1193 => x"00000000",
  1194 => x"52656164",
  1195 => x"696e6720",
  1196 => x"64697265",
  1197 => x"63746f72",
  1198 => x"79207365",
  1199 => x"63746f72",
  1200 => x"2025640a",
  1201 => x"00000000",
  1202 => x"66696c65",
  1203 => x"20222573",
  1204 => x"2220666f",
  1205 => x"756e640d",
  1206 => x"00000000",
  1207 => x"47657446",
  1208 => x"41544c69",
  1209 => x"6e6b2072",
  1210 => x"65747572",
  1211 => x"6e656420",
  1212 => x"25640a00",
  1213 => x"4f70656e",
  1214 => x"65642066",
  1215 => x"696c652c",
  1216 => x"206c6f61",
  1217 => x"64696e67",
  1218 => x"2e2e2e0a",
  1219 => x"00000000",
  1220 => x"52656164",
  1221 => x"696e6720",
  1222 => x"626c6f63",
  1223 => x"6b202564",
  1224 => x"20282564",
  1225 => x"2c202564",
  1226 => x"2c202564",
  1227 => x"292e2e2e",
  1228 => x"00000000",
  1229 => x"626c6f63",
  1230 => x"6b207265",
  1231 => x"61642e0a",
  1232 => x"00000000",
  1233 => x"47657474",
  1234 => x"696e6720",
  1235 => x"6e657874",
  1236 => x"20636c75",
  1237 => x"73746572",
  1238 => x"2e0a0000",
  1239 => x"43616e27",
  1240 => x"74206f70",
  1241 => x"656e2025",
  1242 => x"730a0000",
	others => x"00000000"
);

begin

process (clk)
begin
	if (clk'event and clk = '1') then
		if (from_zpu.memAWriteEnable = '1') and (from_zpu.memBWriteEnable = '1') and (from_zpu.memAAddr=from_zpu.memBAddr) and (from_zpu.memAWrite/=from_zpu.memBWrite) then
			report "write collision" severity failure;
		end if;
	
		if (from_zpu.memAWriteEnable = '1') then
			ram(to_integer(unsigned(from_zpu.memAAddr(maxAddrBitBRAM downto 2)))) := from_zpu.memAWrite;
			to_zpu.memARead <= from_zpu.memAWrite;
		else
			to_zpu.memARead <= ram(to_integer(unsigned(from_zpu.memAAddr(maxAddrBitBRAM downto 2))));
		end if;
	end if;
end process;

process (clk)
begin
	if (clk'event and clk = '1') then
		if (from_zpu.memBWriteEnable = '1') then
			ram(to_integer(unsigned(from_zpu.memBAddr(maxAddrBitBRAM downto 2)))) := from_zpu.memBWrite;
			to_zpu.memBRead <= from_zpu.memBWrite;
		else
			to_zpu.memBRead <= ram(to_integer(unsigned(from_zpu.memBAddr(maxAddrBitBRAM downto 2))));
		end if;
	end if;
end process;


end arch;

