-- ZPU
--
-- Copyright 2004-2008 oharboe - �yvind Harboe - oyvind.harboe@zylin.com
-- Modified by Alastair M. Robinson for the ZPUFlex project.
--
-- The FreeBSD license
-- 
-- Redistribution and use in source and binary forms, with or without
-- modification, are permitted provided that the following conditions
-- are met:
-- 
-- 1. Redistributions of source code must retain the above copyright
--    notice, this list of conditions and the following disclaimer.
-- 2. Redistributions in binary form must reproduce the above
--    copyright notice, this list of conditions and the following
--    disclaimer in the documentation and/or other materials
--    provided with the distribution.
-- 
-- THIS SOFTWARE IS PROVIDED BY THE ZPU PROJECT ``AS IS'' AND ANY
-- EXPRESS OR IMPLIED WARRANTIES, INCLUDING, BUT NOT LIMITED TO,
-- THE IMPLIED WARRANTIES OF MERCHANTABILITY AND FITNESS FOR A
-- PARTICULAR PURPOSE ARE DISCLAIMED. IN NO EVENT SHALL THE
-- ZPU PROJECT OR CONTRIBUTORS BE LIABLE FOR ANY DIRECT,
-- INDIRECT, INCIDENTAL, SPECIAL, EXEMPLARY, OR CONSEQUENTIAL DAMAGES
-- (INCLUDING, BUT NOT LIMITED TO, PROCUREMENT OF SUBSTITUTE GOODS
-- OR SERVICES; LOSS OF USE, DATA, OR PROFITS; OR BUSINESS INTERRUPTION)
-- HOWEVER CAUSED AND ON ANY THEORY OF LIABILITY, WHETHER IN CONTRACT,
-- STRICT LIABILITY, OR TORT (INCLUDING NEGLIGENCE OR OTHERWISE)
-- ARISING IN ANY WAY OUT OF THE USE OF THIS SOFTWARE, EVEN IF
-- ADVISED OF THE POSSIBILITY OF SUCH DAMAGE.
-- 
-- The views and conclusions contained in the software and documentation
-- are those of the authors and should not be interpreted as representing
-- official policies, either expressed or implied, of the ZPU Project.

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;


library work;
use work.zpu_config.all;
use work.zpupkg.all;

entity Interrupt_ROM is
generic
	(
		maxAddrBit : integer := maxAddrBitBRAMLimit -- Specify your actual ROM size to save LEs and unnecessary block RAM usage.
	);
port (
	clk : in std_logic;
	areset : in std_logic := '0';
	from_zpu : in ZPU_ToROM;
	to_zpu : out ZPU_FromROM
);
end Interrupt_ROM;

architecture arch of Interrupt_ROM is

type ram_type is array(natural range 0 to ((2**(maxAddrBit+1))/4)-1) of std_logic_vector(wordSize-1 downto 0);

shared variable ram : ram_type :=
(
     0 => x"0b0b0b88",
     1 => x"dd040000",
     2 => x"00000000",
     3 => x"00000000",
     4 => x"00000000",
     5 => x"00000000",
     6 => x"00000000",
     7 => x"00000000",
     8 => x"88088c08",
     9 => x"90080b0b",
    10 => x"0b88e708",
    11 => x"2d900c8c",
    12 => x"0c880c04",
    13 => x"00000000",
    14 => x"00000000",
    15 => x"00000000",
    16 => x"71fd0608",
    17 => x"72830609",
    18 => x"81058205",
    19 => x"832b2a83",
    20 => x"ffff0652",
    21 => x"04000000",
    22 => x"00000000",
    23 => x"00000000",
    24 => x"71fd0608",
    25 => x"83ffff73",
    26 => x"83060981",
    27 => x"05820583",
    28 => x"2b2b0906",
    29 => x"7383ffff",
    30 => x"0b0b0b0b",
    31 => x"83a50400",
    32 => x"72098105",
    33 => x"72057373",
    34 => x"09060906",
    35 => x"73097306",
    36 => x"070a8106",
    37 => x"53510400",
    38 => x"00000000",
    39 => x"00000000",
    40 => x"72722473",
    41 => x"732e0753",
    42 => x"51040000",
    43 => x"00000000",
    44 => x"00000000",
    45 => x"00000000",
    46 => x"00000000",
    47 => x"00000000",
    48 => x"71737109",
    49 => x"71068106",
    50 => x"09810572",
    51 => x"0a100a72",
    52 => x"0a100a31",
    53 => x"050a8106",
    54 => x"51515351",
    55 => x"04000000",
    56 => x"72722673",
    57 => x"732e0753",
    58 => x"51040000",
    59 => x"00000000",
    60 => x"00000000",
    61 => x"00000000",
    62 => x"00000000",
    63 => x"00000000",
    64 => x"00000000",
    65 => x"00000000",
    66 => x"00000000",
    67 => x"00000000",
    68 => x"00000000",
    69 => x"00000000",
    70 => x"00000000",
    71 => x"00000000",
    72 => x"0b0b0b88",
    73 => x"ba040000",
    74 => x"00000000",
    75 => x"00000000",
    76 => x"00000000",
    77 => x"00000000",
    78 => x"00000000",
    79 => x"00000000",
    80 => x"720a722b",
    81 => x"0a535104",
    82 => x"00000000",
    83 => x"00000000",
    84 => x"00000000",
    85 => x"00000000",
    86 => x"00000000",
    87 => x"00000000",
    88 => x"72729f06",
    89 => x"0981050b",
    90 => x"0b0b889f",
    91 => x"05040000",
    92 => x"00000000",
    93 => x"00000000",
    94 => x"00000000",
    95 => x"00000000",
    96 => x"72722aff",
    97 => x"739f062a",
    98 => x"0974090a",
    99 => x"8106ff05",
   100 => x"06075351",
   101 => x"04000000",
   102 => x"00000000",
   103 => x"00000000",
   104 => x"71715351",
   105 => x"04067383",
   106 => x"06098105",
   107 => x"8205832b",
   108 => x"0b2b0772",
   109 => x"fc060c51",
   110 => x"51040000",
   111 => x"00000000",
   112 => x"72098105",
   113 => x"72050970",
   114 => x"81050906",
   115 => x"0a810653",
   116 => x"51040000",
   117 => x"00000000",
   118 => x"00000000",
   119 => x"00000000",
   120 => x"72098105",
   121 => x"72050970",
   122 => x"81050906",
   123 => x"0a098106",
   124 => x"53510400",
   125 => x"00000000",
   126 => x"00000000",
   127 => x"00000000",
   128 => x"71098105",
   129 => x"52040000",
   130 => x"00000000",
   131 => x"00000000",
   132 => x"00000000",
   133 => x"00000000",
   134 => x"00000000",
   135 => x"00000000",
   136 => x"72720981",
   137 => x"05055351",
   138 => x"04000000",
   139 => x"00000000",
   140 => x"00000000",
   141 => x"00000000",
   142 => x"00000000",
   143 => x"00000000",
   144 => x"72097206",
   145 => x"73730906",
   146 => x"07535104",
   147 => x"00000000",
   148 => x"00000000",
   149 => x"00000000",
   150 => x"00000000",
   151 => x"00000000",
   152 => x"71fc0608",
   153 => x"72830609",
   154 => x"81058305",
   155 => x"1010102a",
   156 => x"81ff0652",
   157 => x"04000000",
   158 => x"00000000",
   159 => x"00000000",
   160 => x"71fc0608",
   161 => x"0b0b0b91",
   162 => x"b4738306",
   163 => x"10100508",
   164 => x"060b0b0b",
   165 => x"88a20400",
   166 => x"00000000",
   167 => x"00000000",
   168 => x"88088c08",
   169 => x"90087575",
   170 => x"0b0b0b8d",
   171 => x"b62d5050",
   172 => x"88085690",
   173 => x"0c8c0c88",
   174 => x"0c510400",
   175 => x"00000000",
   176 => x"88088c08",
   177 => x"90087575",
   178 => x"0b0b0b8e",
   179 => x"e82d5050",
   180 => x"88085690",
   181 => x"0c8c0c88",
   182 => x"0c510400",
   183 => x"00000000",
   184 => x"72097081",
   185 => x"0509060a",
   186 => x"8106ff05",
   187 => x"70547106",
   188 => x"73097274",
   189 => x"05ff0506",
   190 => x"07515151",
   191 => x"04000000",
   192 => x"72097081",
   193 => x"0509060a",
   194 => x"098106ff",
   195 => x"05705471",
   196 => x"06730972",
   197 => x"7405ff05",
   198 => x"06075151",
   199 => x"51040000",
   200 => x"05ff0504",
   201 => x"00000000",
   202 => x"00000000",
   203 => x"00000000",
   204 => x"00000000",
   205 => x"00000000",
   206 => x"00000000",
   207 => x"00000000",
   208 => x"04000000",
   209 => x"00000000",
   210 => x"00000000",
   211 => x"00000000",
   212 => x"00000000",
   213 => x"00000000",
   214 => x"00000000",
   215 => x"00000000",
   216 => x"71810552",
   217 => x"04000000",
   218 => x"00000000",
   219 => x"00000000",
   220 => x"00000000",
   221 => x"00000000",
   222 => x"00000000",
   223 => x"00000000",
   224 => x"00000000",
   225 => x"00000000",
   226 => x"00000000",
   227 => x"00000000",
   228 => x"00000000",
   229 => x"00000000",
   230 => x"00000000",
   231 => x"00000000",
   232 => x"02840572",
   233 => x"10100552",
   234 => x"04000000",
   235 => x"00000000",
   236 => x"00000000",
   237 => x"00000000",
   238 => x"00000000",
   239 => x"00000000",
   240 => x"00000000",
   241 => x"00000000",
   242 => x"00000000",
   243 => x"00000000",
   244 => x"00000000",
   245 => x"00000000",
   246 => x"00000000",
   247 => x"00000000",
   248 => x"717105ff",
   249 => x"05715351",
   250 => x"020d0400",
   251 => x"00000000",
   252 => x"00000000",
   253 => x"00000000",
   254 => x"00000000",
   255 => x"00000000",
   256 => x"10101010",
   257 => x"10101010",
   258 => x"10101010",
   259 => x"10101010",
   260 => x"10101010",
   261 => x"10101010",
   262 => x"10101010",
   263 => x"10101053",
   264 => x"51047381",
   265 => x"ff067383",
   266 => x"06098105",
   267 => x"83051010",
   268 => x"102b0772",
   269 => x"fc060c51",
   270 => x"51047272",
   271 => x"80728106",
   272 => x"ff050972",
   273 => x"06057110",
   274 => x"52720a10",
   275 => x"0a5372ed",
   276 => x"38515153",
   277 => x"51040000",
   278 => x"800488da",
   279 => x"0488da0b",
   280 => x"8cb60404",
   281 => x"00000000",
   282 => x"000463f1",
   283 => x"3d0d923d",
   284 => x"0b0b0b93",
   285 => x"845c5680",
   286 => x"76708405",
   287 => x"5808715f",
   288 => x"5f577d70",
   289 => x"84055f08",
   290 => x"5a805c79",
   291 => x"982a7a88",
   292 => x"2b5b5574",
   293 => x"8638765f",
   294 => x"81f5397c",
   295 => x"802e81cf",
   296 => x"38805d74",
   297 => x"80e42e9b",
   298 => x"387480e4",
   299 => x"268b3874",
   300 => x"80e32e81",
   301 => x"8738818e",
   302 => x"397480f3",
   303 => x"2e80ec38",
   304 => x"81843975",
   305 => x"84177108",
   306 => x"0b0b0b93",
   307 => x"840b0b0b",
   308 => x"0b92b461",
   309 => x"5d585c52",
   310 => x"5753728e",
   311 => x"38b00b0b",
   312 => x"0b0b92b4",
   313 => x"34811454",
   314 => x"ab398a52",
   315 => x"725183a1",
   316 => x"3f880891",
   317 => x"c4053374",
   318 => x"70810556",
   319 => x"348a5272",
   320 => x"5182e93f",
   321 => x"88085388",
   322 => x"08e03873",
   323 => x"0b0b0b92",
   324 => x"b42e9138",
   325 => x"ff145473",
   326 => x"33797081",
   327 => x"055b3481",
   328 => x"1858e839",
   329 => x"80793477",
   330 => x"54ab3975",
   331 => x"84177108",
   332 => x"70545d57",
   333 => x"5380fe3f",
   334 => x"7c549a39",
   335 => x"75841771",
   336 => x"08575753",
   337 => x"b639a551",
   338 => x"80cc3f74",
   339 => x"5180c73f",
   340 => x"821757ae",
   341 => x"3973ff15",
   342 => x"55538073",
   343 => x"25a4387a",
   344 => x"7081055c",
   345 => x"33705255",
   346 => x"ad3f8117",
   347 => x"57e73974",
   348 => x"a52e0981",
   349 => x"06853881",
   350 => x"5d883974",
   351 => x"51983f81",
   352 => x"1757811c",
   353 => x"5c837c25",
   354 => x"fe813874",
   355 => x"fdf4387e",
   356 => x"880c913d",
   357 => x"0d04ff3d",
   358 => x"0d7352c0",
   359 => x"0870882a",
   360 => x"70810651",
   361 => x"51517080",
   362 => x"2ef13871",
   363 => x"c00c7188",
   364 => x"0c833d0d",
   365 => x"04fb3d0d",
   366 => x"77557470",
   367 => x"84055608",
   368 => x"53805472",
   369 => x"982a7388",
   370 => x"2b545271",
   371 => x"802ea238",
   372 => x"c0087088",
   373 => x"2a708106",
   374 => x"51515170",
   375 => x"802ef138",
   376 => x"71c00c81",
   377 => x"16811555",
   378 => x"56837425",
   379 => x"d63871ca",
   380 => x"3875880c",
   381 => x"873d0d04",
   382 => x"7188e70c",
   383 => x"04ffb008",
   384 => x"880c0481",
   385 => x"0bffb00c",
   386 => x"04800bff",
   387 => x"b00c04ff",
   388 => x"3d0df63f",
   389 => x"e83f93c4",
   390 => x"08813270",
   391 => x"93c40c52",
   392 => x"71802e86",
   393 => x"3891d851",
   394 => x"843991e4",
   395 => x"51ff863f",
   396 => x"d23f833d",
   397 => x"0d04803d",
   398 => x"0d800b93",
   399 => x"c40c91f0",
   400 => x"51fef23f",
   401 => x"800bf884",
   402 => x"0c868da0",
   403 => x"0bf8880c",
   404 => x"928851fe",
   405 => x"e03f8c8f",
   406 => x"51ff9d3f",
   407 => x"ffa53f92",
   408 => x"a051fed1",
   409 => x"3f810bf8",
   410 => x"800cff39",
   411 => x"94080294",
   412 => x"0cfd3d0d",
   413 => x"80539408",
   414 => x"8c050852",
   415 => x"94088805",
   416 => x"085182de",
   417 => x"3f880870",
   418 => x"880c5485",
   419 => x"3d0d940c",
   420 => x"04940802",
   421 => x"940cfd3d",
   422 => x"0d815394",
   423 => x"088c0508",
   424 => x"52940888",
   425 => x"05085182",
   426 => x"b93f8808",
   427 => x"70880c54",
   428 => x"853d0d94",
   429 => x"0c049408",
   430 => x"02940cf9",
   431 => x"3d0d800b",
   432 => x"9408fc05",
   433 => x"0c940888",
   434 => x"05088025",
   435 => x"ab389408",
   436 => x"88050830",
   437 => x"94088805",
   438 => x"0c800b94",
   439 => x"08f4050c",
   440 => x"9408fc05",
   441 => x"08883881",
   442 => x"0b9408f4",
   443 => x"050c9408",
   444 => x"f4050894",
   445 => x"08fc050c",
   446 => x"94088c05",
   447 => x"088025ab",
   448 => x"3894088c",
   449 => x"05083094",
   450 => x"088c050c",
   451 => x"800b9408",
   452 => x"f0050c94",
   453 => x"08fc0508",
   454 => x"8838810b",
   455 => x"9408f005",
   456 => x"0c9408f0",
   457 => x"05089408",
   458 => x"fc050c80",
   459 => x"5394088c",
   460 => x"05085294",
   461 => x"08880508",
   462 => x"5181a73f",
   463 => x"88087094",
   464 => x"08f8050c",
   465 => x"549408fc",
   466 => x"0508802e",
   467 => x"8c389408",
   468 => x"f8050830",
   469 => x"9408f805",
   470 => x"0c9408f8",
   471 => x"05087088",
   472 => x"0c54893d",
   473 => x"0d940c04",
   474 => x"94080294",
   475 => x"0cfb3d0d",
   476 => x"800b9408",
   477 => x"fc050c94",
   478 => x"08880508",
   479 => x"80259338",
   480 => x"94088805",
   481 => x"08309408",
   482 => x"88050c81",
   483 => x"0b9408fc",
   484 => x"050c9408",
   485 => x"8c050880",
   486 => x"258c3894",
   487 => x"088c0508",
   488 => x"3094088c",
   489 => x"050c8153",
   490 => x"94088c05",
   491 => x"08529408",
   492 => x"88050851",
   493 => x"ad3f8808",
   494 => x"709408f8",
   495 => x"050c5494",
   496 => x"08fc0508",
   497 => x"802e8c38",
   498 => x"9408f805",
   499 => x"08309408",
   500 => x"f8050c94",
   501 => x"08f80508",
   502 => x"70880c54",
   503 => x"873d0d94",
   504 => x"0c049408",
   505 => x"02940cfd",
   506 => x"3d0d810b",
   507 => x"9408fc05",
   508 => x"0c800b94",
   509 => x"08f8050c",
   510 => x"94088c05",
   511 => x"08940888",
   512 => x"050827ac",
   513 => x"389408fc",
   514 => x"0508802e",
   515 => x"a338800b",
   516 => x"94088c05",
   517 => x"08249938",
   518 => x"94088c05",
   519 => x"08109408",
   520 => x"8c050c94",
   521 => x"08fc0508",
   522 => x"109408fc",
   523 => x"050cc939",
   524 => x"9408fc05",
   525 => x"08802e80",
   526 => x"c9389408",
   527 => x"8c050894",
   528 => x"08880508",
   529 => x"26a13894",
   530 => x"08880508",
   531 => x"94088c05",
   532 => x"08319408",
   533 => x"88050c94",
   534 => x"08f80508",
   535 => x"9408fc05",
   536 => x"08079408",
   537 => x"f8050c94",
   538 => x"08fc0508",
   539 => x"812a9408",
   540 => x"fc050c94",
   541 => x"088c0508",
   542 => x"812a9408",
   543 => x"8c050cff",
   544 => x"af399408",
   545 => x"90050880",
   546 => x"2e8f3894",
   547 => x"08880508",
   548 => x"709408f4",
   549 => x"050c518d",
   550 => x"399408f8",
   551 => x"05087094",
   552 => x"08f4050c",
   553 => x"519408f4",
   554 => x"0508880c",
   555 => x"853d0d94",
   556 => x"0c040000",
   557 => x"00ffffff",
   558 => x"ff00ffff",
   559 => x"ffff00ff",
   560 => x"ffffff00",
   561 => x"30313233",
   562 => x"34353637",
   563 => x"38394142",
   564 => x"43444546",
   565 => x"00000000",
   566 => x"5469636b",
   567 => x"2e2e2e0a",
   568 => x"00000000",
   569 => x"546f636b",
   570 => x"2e2e2e0a",
   571 => x"00000000",
   572 => x"53657474",
   573 => x"696e6720",
   574 => x"75702074",
   575 => x"696d6572",
   576 => x"2e2e2e0a",
   577 => x"00000000",
   578 => x"456e6162",
   579 => x"6c696e67",
   580 => x"20696e74",
   581 => x"65727275",
   582 => x"7074732e",
   583 => x"2e2e0a00",
   584 => x"456e6162",
   585 => x"6c696e67",
   586 => x"2074696d",
   587 => x"65722e2e",
   588 => x"2e0a002e",
	others => x"00000000"
);

begin

process (clk)
begin
	if (clk'event and clk = '1') then
		if (from_zpu.memAWriteEnable = '1') and (from_zpu.memBWriteEnable = '1') and (from_zpu.memAAddr=from_zpu.memBAddr) and (from_zpu.memAWrite/=from_zpu.memBWrite) then
			report "write collision" severity failure;
		end if;
	
		if (from_zpu.memAWriteEnable = '1') then
			ram(to_integer(unsigned(from_zpu.memAAddr(maxAddrBit downto 2)))) := from_zpu.memAWrite;
			to_zpu.memARead <= from_zpu.memAWrite;
		else
			to_zpu.memARead <= ram(to_integer(unsigned(from_zpu.memAAddr(maxAddrBit downto 2))));
		end if;
	end if;
end process;

process (clk)
begin
	if (clk'event and clk = '1') then
		if (from_zpu.memBWriteEnable = '1') then
			ram(to_integer(unsigned(from_zpu.memBAddr(maxAddrBit downto 2)))) := from_zpu.memBWrite;
			to_zpu.memBRead <= from_zpu.memBWrite;
		else
			to_zpu.memBRead <= ram(to_integer(unsigned(from_zpu.memBAddr(maxAddrBit downto 2))));
		end if;
	end if;
end process;


end arch;

