-- ZPU
--
-- Copyright 2004-2008 oharboe - �yvind Harboe - oyvind.harboe@zylin.com
-- Modified by Alastair M. Robinson for the ZPUFlex project.
--
-- The FreeBSD license
-- 
-- Redistribution and use in source and binary forms, with or without
-- modification, are permitted provided that the following conditions
-- are met:
-- 
-- 1. Redistributions of source code must retain the above copyright
--    notice, this list of conditions and the following disclaimer.
-- 2. Redistributions in binary form must reproduce the above
--    copyright notice, this list of conditions and the following
--    disclaimer in the documentation and/or other materials
--    provided with the distribution.
-- 
-- THIS SOFTWARE IS PROVIDED BY THE ZPU PROJECT ``AS IS'' AND ANY
-- EXPRESS OR IMPLIED WARRANTIES, INCLUDING, BUT NOT LIMITED TO,
-- THE IMPLIED WARRANTIES OF MERCHANTABILITY AND FITNESS FOR A
-- PARTICULAR PURPOSE ARE DISCLAIMED. IN NO EVENT SHALL THE
-- ZPU PROJECT OR CONTRIBUTORS BE LIABLE FOR ANY DIRECT,
-- INDIRECT, INCIDENTAL, SPECIAL, EXEMPLARY, OR CONSEQUENTIAL DAMAGES
-- (INCLUDING, BUT NOT LIMITED TO, PROCUREMENT OF SUBSTITUTE GOODS
-- OR SERVICES; LOSS OF USE, DATA, OR PROFITS; OR BUSINESS INTERRUPTION)
-- HOWEVER CAUSED AND ON ANY THEORY OF LIABILITY, WHETHER IN CONTRACT,
-- STRICT LIABILITY, OR TORT (INCLUDING NEGLIGENCE OR OTHERWISE)
-- ARISING IN ANY WAY OUT OF THE USE OF THIS SOFTWARE, EVEN IF
-- ADVISED OF THE POSSIBILITY OF SUCH DAMAGE.
-- 
-- The views and conclusions contained in the software and documentation
-- are those of the authors and should not be interpreted as representing
-- official policies, either expressed or implied, of the ZPU Project.

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;


library work;
use work.zpu_config.all;
use work.zpupkg.all;

entity VGATest_ROM is
generic
	(
		maxAddrBit : integer := maxAddrBitBRAMLimit -- Specify your actual ROM size to save LEs and unnecessary block RAM usage.
	);
port (
	clk : in std_logic;
	areset : in std_logic := '0';
	from_zpu : in ZPU_ToROM;
	to_zpu : out ZPU_FromROM
);
end VGATest_ROM;

architecture arch of VGATest_ROM is

type ram_type is array(natural range 0 to ((2**(maxAddrBit+1))/4)-1) of std_logic_vector(wordSize-1 downto 0);

shared variable ram : ram_type :=
(
     0 => x"0b0b0b88",
     1 => x"dd040000",
     2 => x"00000000",
     3 => x"00000000",
     4 => x"00000000",
     5 => x"00000000",
     6 => x"00000000",
     7 => x"00000000",
     8 => x"04000000",
     9 => x"00000000",
    10 => x"00000000",
    11 => x"00000000",
    12 => x"00000000",
    13 => x"00000000",
    14 => x"00000000",
    15 => x"00000000",
    16 => x"71fd0608",
    17 => x"72830609",
    18 => x"81058205",
    19 => x"832b2a83",
    20 => x"ffff0652",
    21 => x"04000000",
    22 => x"00000000",
    23 => x"00000000",
    24 => x"71fd0608",
    25 => x"83ffff73",
    26 => x"83060981",
    27 => x"05820583",
    28 => x"2b2b0906",
    29 => x"7383ffff",
    30 => x"0b0b0b0b",
    31 => x"83a50400",
    32 => x"72098105",
    33 => x"72057373",
    34 => x"09060906",
    35 => x"73097306",
    36 => x"070a8106",
    37 => x"53510400",
    38 => x"00000000",
    39 => x"00000000",
    40 => x"72722473",
    41 => x"732e0753",
    42 => x"51040000",
    43 => x"00000000",
    44 => x"00000000",
    45 => x"00000000",
    46 => x"00000000",
    47 => x"00000000",
    48 => x"71737109",
    49 => x"71068106",
    50 => x"09810572",
    51 => x"0a100a72",
    52 => x"0a100a31",
    53 => x"050a8106",
    54 => x"51515351",
    55 => x"04000000",
    56 => x"72722673",
    57 => x"732e0753",
    58 => x"51040000",
    59 => x"00000000",
    60 => x"00000000",
    61 => x"00000000",
    62 => x"00000000",
    63 => x"00000000",
    64 => x"00000000",
    65 => x"00000000",
    66 => x"00000000",
    67 => x"00000000",
    68 => x"00000000",
    69 => x"00000000",
    70 => x"00000000",
    71 => x"00000000",
    72 => x"0b0b0b88",
    73 => x"ba040000",
    74 => x"00000000",
    75 => x"00000000",
    76 => x"00000000",
    77 => x"00000000",
    78 => x"00000000",
    79 => x"00000000",
    80 => x"720a722b",
    81 => x"0a535104",
    82 => x"00000000",
    83 => x"00000000",
    84 => x"00000000",
    85 => x"00000000",
    86 => x"00000000",
    87 => x"00000000",
    88 => x"72729f06",
    89 => x"0981050b",
    90 => x"0b0b889f",
    91 => x"05040000",
    92 => x"00000000",
    93 => x"00000000",
    94 => x"00000000",
    95 => x"00000000",
    96 => x"72722aff",
    97 => x"739f062a",
    98 => x"0974090a",
    99 => x"8106ff05",
   100 => x"06075351",
   101 => x"04000000",
   102 => x"00000000",
   103 => x"00000000",
   104 => x"71715351",
   105 => x"04067383",
   106 => x"06098105",
   107 => x"8205832b",
   108 => x"0b2b0772",
   109 => x"fc060c51",
   110 => x"51040000",
   111 => x"00000000",
   112 => x"72098105",
   113 => x"72050970",
   114 => x"81050906",
   115 => x"0a810653",
   116 => x"51040000",
   117 => x"00000000",
   118 => x"00000000",
   119 => x"00000000",
   120 => x"72098105",
   121 => x"72050970",
   122 => x"81050906",
   123 => x"0a098106",
   124 => x"53510400",
   125 => x"00000000",
   126 => x"00000000",
   127 => x"00000000",
   128 => x"71098105",
   129 => x"52040000",
   130 => x"00000000",
   131 => x"00000000",
   132 => x"00000000",
   133 => x"00000000",
   134 => x"00000000",
   135 => x"00000000",
   136 => x"72720981",
   137 => x"05055351",
   138 => x"04000000",
   139 => x"00000000",
   140 => x"00000000",
   141 => x"00000000",
   142 => x"00000000",
   143 => x"00000000",
   144 => x"72097206",
   145 => x"73730906",
   146 => x"07535104",
   147 => x"00000000",
   148 => x"00000000",
   149 => x"00000000",
   150 => x"00000000",
   151 => x"00000000",
   152 => x"71fc0608",
   153 => x"72830609",
   154 => x"81058305",
   155 => x"1010102a",
   156 => x"81ff0652",
   157 => x"04000000",
   158 => x"00000000",
   159 => x"00000000",
   160 => x"71fc0608",
   161 => x"0b0b0b91",
   162 => x"dc738306",
   163 => x"10100508",
   164 => x"060b0b0b",
   165 => x"88a20400",
   166 => x"00000000",
   167 => x"00000000",
   168 => x"88088c08",
   169 => x"90087575",
   170 => x"0b0b0b8d",
   171 => x"de2d5050",
   172 => x"88085690",
   173 => x"0c8c0c88",
   174 => x"0c510400",
   175 => x"00000000",
   176 => x"88088c08",
   177 => x"90087575",
   178 => x"0b0b0b8f",
   179 => x"902d5050",
   180 => x"88085690",
   181 => x"0c8c0c88",
   182 => x"0c510400",
   183 => x"00000000",
   184 => x"72097081",
   185 => x"0509060a",
   186 => x"8106ff05",
   187 => x"70547106",
   188 => x"73097274",
   189 => x"05ff0506",
   190 => x"07515151",
   191 => x"04000000",
   192 => x"72097081",
   193 => x"0509060a",
   194 => x"098106ff",
   195 => x"05705471",
   196 => x"06730972",
   197 => x"7405ff05",
   198 => x"06075151",
   199 => x"51040000",
   200 => x"05ff0504",
   201 => x"00000000",
   202 => x"00000000",
   203 => x"00000000",
   204 => x"00000000",
   205 => x"00000000",
   206 => x"00000000",
   207 => x"00000000",
   208 => x"04000000",
   209 => x"00000000",
   210 => x"00000000",
   211 => x"00000000",
   212 => x"00000000",
   213 => x"00000000",
   214 => x"00000000",
   215 => x"00000000",
   216 => x"71810552",
   217 => x"04000000",
   218 => x"00000000",
   219 => x"00000000",
   220 => x"00000000",
   221 => x"00000000",
   222 => x"00000000",
   223 => x"00000000",
   224 => x"00000000",
   225 => x"00000000",
   226 => x"00000000",
   227 => x"00000000",
   228 => x"00000000",
   229 => x"00000000",
   230 => x"00000000",
   231 => x"00000000",
   232 => x"02840572",
   233 => x"10100552",
   234 => x"04000000",
   235 => x"00000000",
   236 => x"00000000",
   237 => x"00000000",
   238 => x"00000000",
   239 => x"00000000",
   240 => x"00000000",
   241 => x"00000000",
   242 => x"00000000",
   243 => x"00000000",
   244 => x"00000000",
   245 => x"00000000",
   246 => x"00000000",
   247 => x"00000000",
   248 => x"717105ff",
   249 => x"05715351",
   250 => x"020d0400",
   251 => x"00000000",
   252 => x"00000000",
   253 => x"00000000",
   254 => x"00000000",
   255 => x"00000000",
   256 => x"10101010",
   257 => x"10101010",
   258 => x"10101010",
   259 => x"10101010",
   260 => x"10101010",
   261 => x"10101010",
   262 => x"10101010",
   263 => x"10101053",
   264 => x"51047381",
   265 => x"ff067383",
   266 => x"06098105",
   267 => x"83051010",
   268 => x"102b0772",
   269 => x"fc060c51",
   270 => x"51047272",
   271 => x"80728106",
   272 => x"ff050972",
   273 => x"06057110",
   274 => x"52720a10",
   275 => x"0a5372ed",
   276 => x"38515153",
   277 => x"51040000",
   278 => x"800488da",
   279 => x"0488da0b",
   280 => x"8cd20402",
   281 => x"c0050d02",
   282 => x"80c4050b",
   283 => x"0b0b92d0",
   284 => x"5a5c807c",
   285 => x"7084055e",
   286 => x"08715f5f",
   287 => x"577d7084",
   288 => x"055f0856",
   289 => x"80587598",
   290 => x"2a76882b",
   291 => x"57557480",
   292 => x"2e82d038",
   293 => x"7c802eb9",
   294 => x"38805d74",
   295 => x"80e42e81",
   296 => x"9f387480",
   297 => x"e42680dc",
   298 => x"387480e3",
   299 => x"2eba38a5",
   300 => x"518bec2d",
   301 => x"74518bec",
   302 => x"2d821757",
   303 => x"81185883",
   304 => x"7825c338",
   305 => x"74ffb638",
   306 => x"7e880c02",
   307 => x"80c0050d",
   308 => x"0474a52e",
   309 => x"09810698",
   310 => x"38810b81",
   311 => x"19595d83",
   312 => x"7825ffa2",
   313 => x"3889c404",
   314 => x"7b841d71",
   315 => x"08575d5a",
   316 => x"74518bec",
   317 => x"2d811781",
   318 => x"19595783",
   319 => x"7825ff86",
   320 => x"3889c404",
   321 => x"7480f32e",
   322 => x"098106ff",
   323 => x"a2387b84",
   324 => x"1d710870",
   325 => x"545b5d54",
   326 => x"8c8d2d80",
   327 => x"0bff1155",
   328 => x"53807325",
   329 => x"ff963878",
   330 => x"7081055a",
   331 => x"84e02d70",
   332 => x"52558bec",
   333 => x"2d811774",
   334 => x"ff165654",
   335 => x"578aa104",
   336 => x"7b841d71",
   337 => x"080b0b0b",
   338 => x"92d00b0b",
   339 => x"0b0b9280",
   340 => x"615f585e",
   341 => x"525d5372",
   342 => x"ba38b00b",
   343 => x"0b0b0b92",
   344 => x"800b8580",
   345 => x"2d811454",
   346 => x"ff145473",
   347 => x"84e02d7b",
   348 => x"7081055d",
   349 => x"85802d81",
   350 => x"1a5a730b",
   351 => x"0b0b9280",
   352 => x"2e098106",
   353 => x"e338807b",
   354 => x"85802d79",
   355 => x"ff115553",
   356 => x"8aa1048a",
   357 => x"5272518d",
   358 => x"b92d8808",
   359 => x"0b0b0b91",
   360 => x"ec0584e0",
   361 => x"2d747081",
   362 => x"05568580",
   363 => x"2d8a5272",
   364 => x"518d942d",
   365 => x"88085388",
   366 => x"08d93873",
   367 => x"0b0b0b92",
   368 => x"802ec338",
   369 => x"ff145473",
   370 => x"84e02d7b",
   371 => x"7081055d",
   372 => x"85802d81",
   373 => x"1a5a730b",
   374 => x"0b0b9280",
   375 => x"2effa738",
   376 => x"8ae80476",
   377 => x"880c0280",
   378 => x"c0050d04",
   379 => x"02f8050d",
   380 => x"7352c008",
   381 => x"70882a70",
   382 => x"81065151",
   383 => x"5170802e",
   384 => x"f13871c0",
   385 => x"0c71880c",
   386 => x"0288050d",
   387 => x"0402e805",
   388 => x"0d775675",
   389 => x"70840557",
   390 => x"08538054",
   391 => x"72982a73",
   392 => x"882b5452",
   393 => x"71802ea2",
   394 => x"38c00870",
   395 => x"882a7081",
   396 => x"06515151",
   397 => x"70802ef1",
   398 => x"3871c00c",
   399 => x"81158115",
   400 => x"55558374",
   401 => x"25d63871",
   402 => x"ca387488",
   403 => x"0c029805",
   404 => x"0d0402ec",
   405 => x"050d8051",
   406 => x"8480800b",
   407 => x"870a0c81",
   408 => x"11705255",
   409 => x"84808053",
   410 => x"805484fe",
   411 => x"52811170",
   412 => x"83ffff06",
   413 => x"70757084",
   414 => x"05570cfe",
   415 => x"14545151",
   416 => x"718025e9",
   417 => x"38811454",
   418 => x"83df7425",
   419 => x"dd388115",
   420 => x"518cdf04",
   421 => x"94080294",
   422 => x"0cfd3d0d",
   423 => x"80539408",
   424 => x"8c050852",
   425 => x"94088805",
   426 => x"085182de",
   427 => x"3f880870",
   428 => x"880c5485",
   429 => x"3d0d940c",
   430 => x"04940802",
   431 => x"940cfd3d",
   432 => x"0d815394",
   433 => x"088c0508",
   434 => x"52940888",
   435 => x"05085182",
   436 => x"b93f8808",
   437 => x"70880c54",
   438 => x"853d0d94",
   439 => x"0c049408",
   440 => x"02940cf9",
   441 => x"3d0d800b",
   442 => x"9408fc05",
   443 => x"0c940888",
   444 => x"05088025",
   445 => x"ab389408",
   446 => x"88050830",
   447 => x"94088805",
   448 => x"0c800b94",
   449 => x"08f4050c",
   450 => x"9408fc05",
   451 => x"08883881",
   452 => x"0b9408f4",
   453 => x"050c9408",
   454 => x"f4050894",
   455 => x"08fc050c",
   456 => x"94088c05",
   457 => x"088025ab",
   458 => x"3894088c",
   459 => x"05083094",
   460 => x"088c050c",
   461 => x"800b9408",
   462 => x"f0050c94",
   463 => x"08fc0508",
   464 => x"8838810b",
   465 => x"9408f005",
   466 => x"0c9408f0",
   467 => x"05089408",
   468 => x"fc050c80",
   469 => x"5394088c",
   470 => x"05085294",
   471 => x"08880508",
   472 => x"5181a73f",
   473 => x"88087094",
   474 => x"08f8050c",
   475 => x"549408fc",
   476 => x"0508802e",
   477 => x"8c389408",
   478 => x"f8050830",
   479 => x"9408f805",
   480 => x"0c9408f8",
   481 => x"05087088",
   482 => x"0c54893d",
   483 => x"0d940c04",
   484 => x"94080294",
   485 => x"0cfb3d0d",
   486 => x"800b9408",
   487 => x"fc050c94",
   488 => x"08880508",
   489 => x"80259338",
   490 => x"94088805",
   491 => x"08309408",
   492 => x"88050c81",
   493 => x"0b9408fc",
   494 => x"050c9408",
   495 => x"8c050880",
   496 => x"258c3894",
   497 => x"088c0508",
   498 => x"3094088c",
   499 => x"050c8153",
   500 => x"94088c05",
   501 => x"08529408",
   502 => x"88050851",
   503 => x"ad3f8808",
   504 => x"709408f8",
   505 => x"050c5494",
   506 => x"08fc0508",
   507 => x"802e8c38",
   508 => x"9408f805",
   509 => x"08309408",
   510 => x"f8050c94",
   511 => x"08f80508",
   512 => x"70880c54",
   513 => x"873d0d94",
   514 => x"0c049408",
   515 => x"02940cfd",
   516 => x"3d0d810b",
   517 => x"9408fc05",
   518 => x"0c800b94",
   519 => x"08f8050c",
   520 => x"94088c05",
   521 => x"08940888",
   522 => x"050827ac",
   523 => x"389408fc",
   524 => x"0508802e",
   525 => x"a338800b",
   526 => x"94088c05",
   527 => x"08249938",
   528 => x"94088c05",
   529 => x"08109408",
   530 => x"8c050c94",
   531 => x"08fc0508",
   532 => x"109408fc",
   533 => x"050cc939",
   534 => x"9408fc05",
   535 => x"08802e80",
   536 => x"c9389408",
   537 => x"8c050894",
   538 => x"08880508",
   539 => x"26a13894",
   540 => x"08880508",
   541 => x"94088c05",
   542 => x"08319408",
   543 => x"88050c94",
   544 => x"08f80508",
   545 => x"9408fc05",
   546 => x"08079408",
   547 => x"f8050c94",
   548 => x"08fc0508",
   549 => x"812a9408",
   550 => x"fc050c94",
   551 => x"088c0508",
   552 => x"812a9408",
   553 => x"8c050cff",
   554 => x"af399408",
   555 => x"90050880",
   556 => x"2e8f3894",
   557 => x"08880508",
   558 => x"709408f4",
   559 => x"050c518d",
   560 => x"399408f8",
   561 => x"05087094",
   562 => x"08f4050c",
   563 => x"519408f4",
   564 => x"0508880c",
   565 => x"853d0d94",
   566 => x"0c040000",
   567 => x"00ffffff",
   568 => x"ff00ffff",
   569 => x"ffff00ff",
   570 => x"ffffff00",
   571 => x"30313233",
   572 => x"34353637",
   573 => x"38394142",
   574 => x"43444546",
   575 => x"00000000",
	others => x"00000000"
);

begin

process (clk)
begin
	if (clk'event and clk = '1') then
		if (from_zpu.memAWriteEnable = '1') and (from_zpu.memBWriteEnable = '1') and (from_zpu.memAAddr=from_zpu.memBAddr) and (from_zpu.memAWrite/=from_zpu.memBWrite) then
			report "write collision" severity failure;
		end if;
	
		if (from_zpu.memAWriteEnable = '1') then
			ram(to_integer(unsigned(from_zpu.memAAddr(maxAddrBit downto 2)))) := from_zpu.memAWrite;
			to_zpu.memARead <= from_zpu.memAWrite;
		else
			to_zpu.memARead <= ram(to_integer(unsigned(from_zpu.memAAddr(maxAddrBit downto 2))));
		end if;
	end if;
end process;

process (clk)
begin
	if (clk'event and clk = '1') then
		if (from_zpu.memBWriteEnable = '1') then
			ram(to_integer(unsigned(from_zpu.memBAddr(maxAddrBit downto 2)))) := from_zpu.memBWrite;
			to_zpu.memBRead <= from_zpu.memBWrite;
		else
			to_zpu.memBRead <= ram(to_integer(unsigned(from_zpu.memBAddr(maxAddrBit downto 2))));
		end if;
	end if;
end process;


end arch;

