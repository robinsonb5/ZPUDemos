-- ZPU
--
-- Copyright 2004-2008 oharboe - �yvind Harboe - oyvind.harboe@zylin.com
-- Modified by Alastair M. Robinson for the ZPUFlex project.
--
-- The FreeBSD license
-- 
-- Redistribution and use in source and binary forms, with or without
-- modification, are permitted provided that the following conditions
-- are met:
-- 
-- 1. Redistributions of source code must retain the above copyright
--    notice, this list of conditions and the following disclaimer.
-- 2. Redistributions in binary form must reproduce the above
--    copyright notice, this list of conditions and the following
--    disclaimer in the documentation and/or other materials
--    provided with the distribution.
-- 
-- THIS SOFTWARE IS PROVIDED BY THE ZPU PROJECT ``AS IS'' AND ANY
-- EXPRESS OR IMPLIED WARRANTIES, INCLUDING, BUT NOT LIMITED TO,
-- THE IMPLIED WARRANTIES OF MERCHANTABILITY AND FITNESS FOR A
-- PARTICULAR PURPOSE ARE DISCLAIMED. IN NO EVENT SHALL THE
-- ZPU PROJECT OR CONTRIBUTORS BE LIABLE FOR ANY DIRECT,
-- INDIRECT, INCIDENTAL, SPECIAL, EXEMPLARY, OR CONSEQUENTIAL DAMAGES
-- (INCLUDING, BUT NOT LIMITED TO, PROCUREMENT OF SUBSTITUTE GOODS
-- OR SERVICES; LOSS OF USE, DATA, OR PROFITS; OR BUSINESS INTERRUPTION)
-- HOWEVER CAUSED AND ON ANY THEORY OF LIABILITY, WHETHER IN CONTRACT,
-- STRICT LIABILITY, OR TORT (INCLUDING NEGLIGENCE OR OTHERWISE)
-- ARISING IN ANY WAY OUT OF THE USE OF THIS SOFTWARE, EVEN IF
-- ADVISED OF THE POSSIBILITY OF SUCH DAMAGE.
-- 
-- The views and conclusions contained in the software and documentation
-- are those of the authors and should not be interpreted as representing
-- official policies, either expressed or implied, of the ZPU Project.

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;


library work;
use work.zpupkg.all;

entity SDBootstrap_ROM is
generic
	(
		maxAddrBitBRAM : integer := maxAddrBitBRAMLimit -- Specify your actual ROM size to save LEs and unnecessary block RAM usage.
	);
port (
	clk : in std_logic;
	areset : in std_logic := '0';
	from_zpu : in ZPU_ToROM;
	to_zpu : out ZPU_FromROM
);
end SDBootstrap_ROM;

architecture arch of SDBootstrap_ROM is

type ram_type is array(natural range 0 to ((2**(maxAddrBitBRAM+1))/4)-1) of std_logic_vector(wordSize-1 downto 0);

shared variable ram : ram_type :=
(
     0 => x"84808080",
     1 => x"8c0b8480",
     2 => x"8081e004",
     3 => x"00848080",
     4 => x"808c04ff",
     5 => x"0d800404",
     6 => x"40000017",
     7 => x"00000000",
     8 => x"0b83ffe0",
     9 => x"80080b83",
    10 => x"ffe08408",
    11 => x"0b83ffe0",
    12 => x"88088480",
    13 => x"80809808",
    14 => x"2d0b83ff",
    15 => x"e0880c0b",
    16 => x"83ffe084",
    17 => x"0c0b83ff",
    18 => x"e0800c04",
    19 => x"00000000",
    20 => x"00000000",
    21 => x"00000000",
    22 => x"00000000",
    23 => x"00000000",
    24 => x"71fd0608",
    25 => x"72830609",
    26 => x"81058205",
    27 => x"832b2a83",
    28 => x"ffff0652",
    29 => x"0471fc06",
    30 => x"08728306",
    31 => x"09810583",
    32 => x"05101010",
    33 => x"2a81ff06",
    34 => x"520471fd",
    35 => x"060883ff",
    36 => x"ff738306",
    37 => x"09810582",
    38 => x"05832b2b",
    39 => x"09067383",
    40 => x"ffff0673",
    41 => x"83060981",
    42 => x"05820583",
    43 => x"2b0b2b07",
    44 => x"72fc060c",
    45 => x"51510471",
    46 => x"fc060884",
    47 => x"8080a1cc",
    48 => x"73830610",
    49 => x"10050806",
    50 => x"7381ff06",
    51 => x"73830609",
    52 => x"81058305",
    53 => x"1010102b",
    54 => x"0772fc06",
    55 => x"0c515104",
    56 => x"83ffe080",
    57 => x"7083fff5",
    58 => x"f0278e38",
    59 => x"80717084",
    60 => x"05530c84",
    61 => x"808081e4",
    62 => x"04848080",
    63 => x"808c5184",
    64 => x"80808fc7",
    65 => x"0402ec05",
    66 => x"0d765380",
    67 => x"5572752e",
    68 => x"be388754",
    69 => x"729c2a73",
    70 => x"842b5452",
    71 => x"71802e83",
    72 => x"38815589",
    73 => x"72258a38",
    74 => x"b7125284",
    75 => x"808082b4",
    76 => x"04b01252",
    77 => x"74802e89",
    78 => x"38715184",
    79 => x"808085a1",
    80 => x"2dff1454",
    81 => x"738025cc",
    82 => x"38848080",
    83 => x"82d704b0",
    84 => x"51848080",
    85 => x"85a12d80",
    86 => x"0b83ffe0",
    87 => x"800c0294",
    88 => x"050d0402",
    89 => x"c0050d02",
    90 => x"80c40557",
    91 => x"80707870",
    92 => x"84055a08",
    93 => x"72415f5d",
    94 => x"587c7084",
    95 => x"055e085a",
    96 => x"805b7998",
    97 => x"2a7a882b",
    98 => x"5b567589",
    99 => x"38775f84",
   100 => x"80808595",
   101 => x"047d802e",
   102 => x"81d33880",
   103 => x"5e7580e4",
   104 => x"2e8a3875",
   105 => x"80f82e09",
   106 => x"81068938",
   107 => x"76841871",
   108 => x"085e5854",
   109 => x"7580e42e",
   110 => x"a6387580",
   111 => x"e4268e38",
   112 => x"7580e32e",
   113 => x"80d93884",
   114 => x"808084ad",
   115 => x"047580f3",
   116 => x"2eb53875",
   117 => x"80f82e8f",
   118 => x"38848080",
   119 => x"84ad048a",
   120 => x"53848080",
   121 => x"83e90490",
   122 => x"5383ffe0",
   123 => x"e0527b51",
   124 => x"84808082",
   125 => x"852d83ff",
   126 => x"e0800883",
   127 => x"ffe0e05a",
   128 => x"55848080",
   129 => x"84c60476",
   130 => x"84187108",
   131 => x"70545b58",
   132 => x"54848080",
   133 => x"85c52d80",
   134 => x"55848080",
   135 => x"84c60476",
   136 => x"84187108",
   137 => x"58585484",
   138 => x"808084fd",
   139 => x"04a55184",
   140 => x"808085a1",
   141 => x"2d755184",
   142 => x"808085a1",
   143 => x"2d821858",
   144 => x"84808085",
   145 => x"880474ff",
   146 => x"16565480",
   147 => x"7425b938",
   148 => x"78708105",
   149 => x"5a848080",
   150 => x"80f52d70",
   151 => x"52568480",
   152 => x"8085a12d",
   153 => x"81185884",
   154 => x"808084c6",
   155 => x"0475a52e",
   156 => x"09810689",
   157 => x"38815e84",
   158 => x"80808588",
   159 => x"04755184",
   160 => x"808085a1",
   161 => x"2d811858",
   162 => x"811b5b83",
   163 => x"7b25fdf2",
   164 => x"3875fde5",
   165 => x"387e83ff",
   166 => x"e0800c02",
   167 => x"80c0050d",
   168 => x"0402f805",
   169 => x"0d7352c0",
   170 => x"0870882a",
   171 => x"70810651",
   172 => x"51517080",
   173 => x"2ef13871",
   174 => x"c00c7183",
   175 => x"ffe0800c",
   176 => x"0288050d",
   177 => x"0402e805",
   178 => x"0d807857",
   179 => x"55757084",
   180 => x"05570853",
   181 => x"80547298",
   182 => x"2a73882b",
   183 => x"54527180",
   184 => x"2ea238c0",
   185 => x"0870882a",
   186 => x"70810651",
   187 => x"51517080",
   188 => x"2ef13871",
   189 => x"c00c8115",
   190 => x"81155555",
   191 => x"837425d6",
   192 => x"3871ca38",
   193 => x"7483ffe0",
   194 => x"800c0298",
   195 => x"050d0402",
   196 => x"f4050dd4",
   197 => x"5281ff72",
   198 => x"0c710853",
   199 => x"81ff720c",
   200 => x"72882b83",
   201 => x"fe800672",
   202 => x"087081ff",
   203 => x"06515253",
   204 => x"81ff720c",
   205 => x"72710788",
   206 => x"2b720870",
   207 => x"81ff0651",
   208 => x"525381ff",
   209 => x"720c7271",
   210 => x"07882b72",
   211 => x"087081ff",
   212 => x"06720783",
   213 => x"ffe0800c",
   214 => x"5253028c",
   215 => x"050d0402",
   216 => x"f4050d74",
   217 => x"767181ff",
   218 => x"06d40c53",
   219 => x"5383fff1",
   220 => x"a0088538",
   221 => x"71892b52",
   222 => x"71982ad4",
   223 => x"0c71902a",
   224 => x"7081ff06",
   225 => x"d40c5171",
   226 => x"882a7081",
   227 => x"ff06d40c",
   228 => x"517181ff",
   229 => x"06d40c72",
   230 => x"902a7081",
   231 => x"ff06d40c",
   232 => x"51d40870",
   233 => x"81ff0651",
   234 => x"5182b8bf",
   235 => x"527081ff",
   236 => x"2e098106",
   237 => x"943881ff",
   238 => x"0bd40cd4",
   239 => x"087081ff",
   240 => x"06ff1454",
   241 => x"515171e5",
   242 => x"387083ff",
   243 => x"e0800c02",
   244 => x"8c050d04",
   245 => x"02fc050d",
   246 => x"81c75181",
   247 => x"ff0bd40c",
   248 => x"ff115170",
   249 => x"8025f438",
   250 => x"0284050d",
   251 => x"0402f005",
   252 => x"0d848080",
   253 => x"87d42d81",
   254 => x"9c9f5380",
   255 => x"5287fc80",
   256 => x"f7518480",
   257 => x"8086df2d",
   258 => x"83ffe080",
   259 => x"085483ff",
   260 => x"e0800881",
   261 => x"2e098106",
   262 => x"ae3881ff",
   263 => x"0bd40c82",
   264 => x"0a52849c",
   265 => x"80e95184",
   266 => x"808086df",
   267 => x"2d83ffe0",
   268 => x"80088e38",
   269 => x"81ff0bd4",
   270 => x"0c735384",
   271 => x"808088ce",
   272 => x"04848080",
   273 => x"87d42dff",
   274 => x"135372ff",
   275 => x"ae387283",
   276 => x"ffe0800c",
   277 => x"0290050d",
   278 => x"0402f405",
   279 => x"0d81ff0b",
   280 => x"d40c8480",
   281 => x"80a1dc51",
   282 => x"84808085",
   283 => x"c52d9353",
   284 => x"805287fc",
   285 => x"80c15184",
   286 => x"808086df",
   287 => x"2d83ffe0",
   288 => x"80088e38",
   289 => x"81ff0bd4",
   290 => x"0c815384",
   291 => x"8080899d",
   292 => x"04848080",
   293 => x"87d42dff",
   294 => x"135372d4",
   295 => x"387283ff",
   296 => x"e0800c02",
   297 => x"8c050d04",
   298 => x"02f0050d",
   299 => x"84808087",
   300 => x"d42d83aa",
   301 => x"52849c80",
   302 => x"c8518480",
   303 => x"8086df2d",
   304 => x"83ffe080",
   305 => x"0883ffe0",
   306 => x"80085384",
   307 => x"8080a1e8",
   308 => x"52538480",
   309 => x"8082e32d",
   310 => x"72812e09",
   311 => x"8106a938",
   312 => x"84808086",
   313 => x"8f2d83ff",
   314 => x"e0800883",
   315 => x"ffff0653",
   316 => x"7283aa2e",
   317 => x"bb3883ff",
   318 => x"e0800852",
   319 => x"848080a2",
   320 => x"80518480",
   321 => x"8082e32d",
   322 => x"84808088",
   323 => x"d92d8480",
   324 => x"808aa804",
   325 => x"81548480",
   326 => x"808bd304",
   327 => x"848080a2",
   328 => x"98518480",
   329 => x"8082e32d",
   330 => x"80548480",
   331 => x"808bd304",
   332 => x"81ff0bd4",
   333 => x"0cb15384",
   334 => x"808087ed",
   335 => x"2d83ffe0",
   336 => x"8008802e",
   337 => x"80fe3880",
   338 => x"5287fc80",
   339 => x"fa518480",
   340 => x"8086df2d",
   341 => x"83ffe080",
   342 => x"0880d738",
   343 => x"83ffe080",
   344 => x"08528480",
   345 => x"80a2b451",
   346 => x"84808082",
   347 => x"e32d81ff",
   348 => x"0bd40cd4",
   349 => x"087081ff",
   350 => x"06705484",
   351 => x"8080a2c0",
   352 => x"53515384",
   353 => x"808082e3",
   354 => x"2d81ff0b",
   355 => x"d40c81ff",
   356 => x"0bd40c81",
   357 => x"ff0bd40c",
   358 => x"81ff0bd4",
   359 => x"0c72862a",
   360 => x"70810670",
   361 => x"56515372",
   362 => x"802ea838",
   363 => x"8480808a",
   364 => x"940483ff",
   365 => x"e0800852",
   366 => x"848080a2",
   367 => x"b4518480",
   368 => x"8082e32d",
   369 => x"72822efe",
   370 => x"d338ff13",
   371 => x"5372fee7",
   372 => x"38725473",
   373 => x"83ffe080",
   374 => x"0c029005",
   375 => x"0d0402f4",
   376 => x"050d810b",
   377 => x"83fff1a0",
   378 => x"0cd00870",
   379 => x"8f2a7081",
   380 => x"06515153",
   381 => x"72f33872",
   382 => x"d00c8480",
   383 => x"8087d42d",
   384 => x"848080a2",
   385 => x"d0518480",
   386 => x"8085c52d",
   387 => x"d008708f",
   388 => x"2a708106",
   389 => x"51515372",
   390 => x"f338810b",
   391 => x"d00c8753",
   392 => x"805284d4",
   393 => x"80c05184",
   394 => x"808086df",
   395 => x"2d83ffe0",
   396 => x"8008812e",
   397 => x"97387282",
   398 => x"2e098106",
   399 => x"89388053",
   400 => x"8480808d",
   401 => x"8d04ff13",
   402 => x"5372d538",
   403 => x"84808089",
   404 => x"a82d83ff",
   405 => x"e0800883",
   406 => x"fff1a00c",
   407 => x"83ffe080",
   408 => x"088e3881",
   409 => x"5287fc80",
   410 => x"d0518480",
   411 => x"8086df2d",
   412 => x"81ff0bd4",
   413 => x"0cd00870",
   414 => x"8f2a7081",
   415 => x"06515153",
   416 => x"72f33872",
   417 => x"d00c81ff",
   418 => x"0bd40c81",
   419 => x"537283ff",
   420 => x"e0800c02",
   421 => x"8c050d04",
   422 => x"800b83ff",
   423 => x"e0800c04",
   424 => x"02e0050d",
   425 => x"797b5757",
   426 => x"805881ff",
   427 => x"0bd40cd0",
   428 => x"08708f2a",
   429 => x"70810651",
   430 => x"515473f3",
   431 => x"3882810b",
   432 => x"d00c81ff",
   433 => x"0bd40c76",
   434 => x"5287fc80",
   435 => x"d1518480",
   436 => x"8086df2d",
   437 => x"80dbc6df",
   438 => x"5583ffe0",
   439 => x"8008802e",
   440 => x"9b3883ff",
   441 => x"e0800853",
   442 => x"76528480",
   443 => x"80a2dc51",
   444 => x"84808082",
   445 => x"e32d8480",
   446 => x"808ed204",
   447 => x"81ff0bd4",
   448 => x"0cd40870",
   449 => x"81ff0651",
   450 => x"547381fe",
   451 => x"2e098106",
   452 => x"a53880ff",
   453 => x"54848080",
   454 => x"868f2d83",
   455 => x"ffe08008",
   456 => x"76708405",
   457 => x"580cff14",
   458 => x"54738025",
   459 => x"e8388158",
   460 => x"8480808e",
   461 => x"bc04ff15",
   462 => x"5574c138",
   463 => x"81ff0bd4",
   464 => x"0cd00870",
   465 => x"8f2a7081",
   466 => x"06515154",
   467 => x"73f33873",
   468 => x"d00c7783",
   469 => x"ffe0800c",
   470 => x"02a0050d",
   471 => x"0402f405",
   472 => x"0d747088",
   473 => x"2a83fe80",
   474 => x"06707298",
   475 => x"2a077288",
   476 => x"2b87fc80",
   477 => x"80067398",
   478 => x"2b81f00a",
   479 => x"06717307",
   480 => x"0783ffe0",
   481 => x"800c5651",
   482 => x"5351028c",
   483 => x"050d0402",
   484 => x"f8050d02",
   485 => x"8e058480",
   486 => x"8080f52d",
   487 => x"74882b07",
   488 => x"7083ffff",
   489 => x"0683ffe0",
   490 => x"800c5102",
   491 => x"88050d04",
   492 => x"02f8050d",
   493 => x"7370902b",
   494 => x"71902a07",
   495 => x"83ffe080",
   496 => x"0c520288",
   497 => x"050d0402",
   498 => x"ec050d80",
   499 => x"0bfc800c",
   500 => x"848080a2",
   501 => x"fc518480",
   502 => x"8085c52d",
   503 => x"8480808b",
   504 => x"de2d83ff",
   505 => x"e0800880",
   506 => x"2e828638",
   507 => x"848080a3",
   508 => x"94518480",
   509 => x"8085c52d",
   510 => x"84808092",
   511 => x"d52d83ff",
   512 => x"e1a05284",
   513 => x"8080a3ac",
   514 => x"51848080",
   515 => x"a0a82d83",
   516 => x"ffe08008",
   517 => x"802e81cd",
   518 => x"3883ffe1",
   519 => x"a00b8480",
   520 => x"80a3b852",
   521 => x"54848080",
   522 => x"85c52d80",
   523 => x"55737081",
   524 => x"05558480",
   525 => x"8080f52d",
   526 => x"5372a02e",
   527 => x"80e63872",
   528 => x"c00c72a3",
   529 => x"2e818438",
   530 => x"7280c72e",
   531 => x"0981068d",
   532 => x"38848080",
   533 => x"80932d84",
   534 => x"808090ff",
   535 => x"04728a2e",
   536 => x"0981068d",
   537 => x"38848080",
   538 => x"808c2d84",
   539 => x"808090ff",
   540 => x"047280cc",
   541 => x"2e098106",
   542 => x"863883ff",
   543 => x"e1a05472",
   544 => x"81df06f0",
   545 => x"057081ff",
   546 => x"065153b8",
   547 => x"73278938",
   548 => x"ef137081",
   549 => x"ff065153",
   550 => x"74842b73",
   551 => x"07558480",
   552 => x"8090ad04",
   553 => x"72a32ea3",
   554 => x"38737081",
   555 => x"05558480",
   556 => x"8080f52d",
   557 => x"5372a02e",
   558 => x"f038ff14",
   559 => x"75537052",
   560 => x"54848080",
   561 => x"a0a82d74",
   562 => x"fc800c73",
   563 => x"70810555",
   564 => x"84808080",
   565 => x"f52d5372",
   566 => x"8a2e0981",
   567 => x"06ed3884",
   568 => x"808090ab",
   569 => x"04848080",
   570 => x"a3cc5184",
   571 => x"808085c5",
   572 => x"2d848080",
   573 => x"a3e85184",
   574 => x"808085c5",
   575 => x"2d800b83",
   576 => x"ffe0800c",
   577 => x"0294050d",
   578 => x"0402e805",
   579 => x"0d77797b",
   580 => x"58555580",
   581 => x"53727625",
   582 => x"af387470",
   583 => x"81055684",
   584 => x"808080f5",
   585 => x"2d747081",
   586 => x"05568480",
   587 => x"8080f52d",
   588 => x"52527171",
   589 => x"2e893881",
   590 => x"51848080",
   591 => x"92ca0481",
   592 => x"13538480",
   593 => x"80929504",
   594 => x"80517083",
   595 => x"ffe0800c",
   596 => x"0298050d",
   597 => x"0402d805",
   598 => x"0d800b83",
   599 => x"fff5dc0c",
   600 => x"848080a3",
   601 => x"f4518480",
   602 => x"8085c52d",
   603 => x"83fff1b8",
   604 => x"52805184",
   605 => x"80808da0",
   606 => x"2d83ffe0",
   607 => x"80085483",
   608 => x"ffe08008",
   609 => x"95388480",
   610 => x"80a48451",
   611 => x"84808085",
   612 => x"c52d7355",
   613 => x"8480809b",
   614 => x"84048480",
   615 => x"80a49851",
   616 => x"84808085",
   617 => x"c52d8056",
   618 => x"810b83ff",
   619 => x"f1ac0c88",
   620 => x"53848080",
   621 => x"a4b05283",
   622 => x"fff1ee51",
   623 => x"84808092",
   624 => x"892d83ff",
   625 => x"e0800876",
   626 => x"2e098106",
   627 => x"8b3883ff",
   628 => x"e0800883",
   629 => x"fff1ac0c",
   630 => x"88538480",
   631 => x"80a4bc52",
   632 => x"83fff28a",
   633 => x"51848080",
   634 => x"92892d83",
   635 => x"ffe08008",
   636 => x"8b3883ff",
   637 => x"e0800883",
   638 => x"fff1ac0c",
   639 => x"83fff1ac",
   640 => x"08528480",
   641 => x"80a4c851",
   642 => x"84808082",
   643 => x"e32d83ff",
   644 => x"f1ac0880",
   645 => x"2e81cb38",
   646 => x"83fff4fe",
   647 => x"0b848080",
   648 => x"80f52d83",
   649 => x"fff4ff0b",
   650 => x"84808080",
   651 => x"f52d7198",
   652 => x"2b71902b",
   653 => x"0783fff5",
   654 => x"800b8480",
   655 => x"8080f52d",
   656 => x"70882b72",
   657 => x"0783fff5",
   658 => x"810b8480",
   659 => x"8080f52d",
   660 => x"710783ff",
   661 => x"f5b60b84",
   662 => x"808080f5",
   663 => x"2d83fff5",
   664 => x"b70b8480",
   665 => x"8080f52d",
   666 => x"71882b07",
   667 => x"535f5452",
   668 => x"5a565755",
   669 => x"7381abaa",
   670 => x"2e098106",
   671 => x"95387551",
   672 => x"8480808e",
   673 => x"dd2d83ff",
   674 => x"e0800856",
   675 => x"84808095",
   676 => x"ab047382",
   677 => x"d4d52e93",
   678 => x"38848080",
   679 => x"a4dc5184",
   680 => x"808085c5",
   681 => x"2d848080",
   682 => x"97b70475",
   683 => x"52848080",
   684 => x"a4fc5184",
   685 => x"808082e3",
   686 => x"2d83fff1",
   687 => x"b8527551",
   688 => x"8480808d",
   689 => x"a02d83ff",
   690 => x"e0800855",
   691 => x"83ffe080",
   692 => x"08802e85",
   693 => x"af388480",
   694 => x"80a59451",
   695 => x"84808085",
   696 => x"c52d8480",
   697 => x"80a5bc51",
   698 => x"84808082",
   699 => x"e32d8853",
   700 => x"848080a4",
   701 => x"bc5283ff",
   702 => x"f28a5184",
   703 => x"80809289",
   704 => x"2d83ffe0",
   705 => x"80088e38",
   706 => x"810b83ff",
   707 => x"f5dc0c84",
   708 => x"808096c3",
   709 => x"04885384",
   710 => x"8080a4b0",
   711 => x"5283fff1",
   712 => x"ee518480",
   713 => x"8092892d",
   714 => x"83ffe080",
   715 => x"08802e93",
   716 => x"38848080",
   717 => x"a5d45184",
   718 => x"808082e3",
   719 => x"2d848080",
   720 => x"97b70483",
   721 => x"fff5b60b",
   722 => x"84808080",
   723 => x"f52d5473",
   724 => x"80d52e09",
   725 => x"810680df",
   726 => x"3883fff5",
   727 => x"b70b8480",
   728 => x"8080f52d",
   729 => x"547381aa",
   730 => x"2e098106",
   731 => x"80c93880",
   732 => x"0b83fff1",
   733 => x"b80b8480",
   734 => x"8080f52d",
   735 => x"56547481",
   736 => x"e92e8338",
   737 => x"81547481",
   738 => x"eb2e8c38",
   739 => x"80557375",
   740 => x"2e098106",
   741 => x"83ee3883",
   742 => x"fff1c30b",
   743 => x"84808080",
   744 => x"f52d5978",
   745 => x"923883ff",
   746 => x"f1c40b84",
   747 => x"808080f5",
   748 => x"2d547382",
   749 => x"2e893880",
   750 => x"55848080",
   751 => x"9b840483",
   752 => x"fff1c50b",
   753 => x"84808080",
   754 => x"f52d7083",
   755 => x"fff5e40c",
   756 => x"ff117083",
   757 => x"fff5d80c",
   758 => x"54528480",
   759 => x"80a5f451",
   760 => x"84808082",
   761 => x"e32d83ff",
   762 => x"f1c60b84",
   763 => x"808080f5",
   764 => x"2d83fff1",
   765 => x"c70b8480",
   766 => x"8080f52d",
   767 => x"56760575",
   768 => x"82802905",
   769 => x"7083fff5",
   770 => x"cc0c83ff",
   771 => x"f1c80b84",
   772 => x"808080f5",
   773 => x"2d7083ff",
   774 => x"f5c80c83",
   775 => x"fff5dc08",
   776 => x"59575876",
   777 => x"802e81ec",
   778 => x"38885384",
   779 => x"8080a4bc",
   780 => x"5283fff2",
   781 => x"8a518480",
   782 => x"8092892d",
   783 => x"785583ff",
   784 => x"e0800882",
   785 => x"bf3883ff",
   786 => x"f5e40870",
   787 => x"842b83ff",
   788 => x"f5b80c70",
   789 => x"83fff5e0",
   790 => x"0c83fff1",
   791 => x"dd0b8480",
   792 => x"8080f52d",
   793 => x"83fff1dc",
   794 => x"0b848080",
   795 => x"80f52d71",
   796 => x"82802905",
   797 => x"83fff1de",
   798 => x"0b848080",
   799 => x"80f52d70",
   800 => x"84808029",
   801 => x"1283fff1",
   802 => x"df0b8480",
   803 => x"8080f52d",
   804 => x"7081800a",
   805 => x"29127083",
   806 => x"fff1b00c",
   807 => x"83fff5c8",
   808 => x"08712983",
   809 => x"fff5cc08",
   810 => x"057083ff",
   811 => x"f5ec0c83",
   812 => x"fff1e50b",
   813 => x"84808080",
   814 => x"f52d83ff",
   815 => x"f1e40b84",
   816 => x"808080f5",
   817 => x"2d718280",
   818 => x"290583ff",
   819 => x"f1e60b84",
   820 => x"808080f5",
   821 => x"2d708480",
   822 => x"80291283",
   823 => x"fff1e70b",
   824 => x"84808080",
   825 => x"f52d7098",
   826 => x"2b81f00a",
   827 => x"06720570",
   828 => x"83fff1b4",
   829 => x"0cfe117e",
   830 => x"29770583",
   831 => x"fff5d40c",
   832 => x"52575257",
   833 => x"5d575152",
   834 => x"5f525c57",
   835 => x"57578480",
   836 => x"809b8204",
   837 => x"83fff1ca",
   838 => x"0b848080",
   839 => x"80f52d83",
   840 => x"fff1c90b",
   841 => x"84808080",
   842 => x"f52d7182",
   843 => x"80290570",
   844 => x"83fff5b8",
   845 => x"0c70a029",
   846 => x"83ff0570",
   847 => x"892a7083",
   848 => x"fff5e00c",
   849 => x"83fff1cf",
   850 => x"0b848080",
   851 => x"80f52d83",
   852 => x"fff1ce0b",
   853 => x"84808080",
   854 => x"f52d7182",
   855 => x"80290570",
   856 => x"83fff1b0",
   857 => x"0c7b7129",
   858 => x"1e7083ff",
   859 => x"f5d40c7d",
   860 => x"83fff1b4",
   861 => x"0c730583",
   862 => x"fff5ec0c",
   863 => x"555e5151",
   864 => x"55558155",
   865 => x"7483ffe0",
   866 => x"800c02a8",
   867 => x"050d0402",
   868 => x"ec050d76",
   869 => x"70872c71",
   870 => x"80ff0657",
   871 => x"555383ff",
   872 => x"f5dc088a",
   873 => x"3872882c",
   874 => x"7381ff06",
   875 => x"565483ff",
   876 => x"f5cc0814",
   877 => x"52848080",
   878 => x"a6985184",
   879 => x"808082e3",
   880 => x"2d83fff1",
   881 => x"b85283ff",
   882 => x"f5cc0814",
   883 => x"51848080",
   884 => x"8da02d83",
   885 => x"ffe08008",
   886 => x"5383ffe0",
   887 => x"8008802e",
   888 => x"80c93883",
   889 => x"fff5dc08",
   890 => x"802ea238",
   891 => x"74842983",
   892 => x"fff1b805",
   893 => x"70085253",
   894 => x"8480808e",
   895 => x"dd2d83ff",
   896 => x"e08008f0",
   897 => x"0a065584",
   898 => x"80809ca9",
   899 => x"04741083",
   900 => x"fff1b805",
   901 => x"70848080",
   902 => x"80e02d52",
   903 => x"53848080",
   904 => x"8f8f2d83",
   905 => x"ffe08008",
   906 => x"55745372",
   907 => x"83ffe080",
   908 => x"0c029405",
   909 => x"0d0402c8",
   910 => x"050d7f61",
   911 => x"5f5c800b",
   912 => x"83fff1b4",
   913 => x"0883fff5",
   914 => x"d4085859",
   915 => x"5783fff5",
   916 => x"dc08772e",
   917 => x"8f3883ff",
   918 => x"f5e40884",
   919 => x"2b598480",
   920 => x"809cec04",
   921 => x"83fff5e0",
   922 => x"08842b59",
   923 => x"805a7979",
   924 => x"2781dc38",
   925 => x"798f06a0",
   926 => x"18585473",
   927 => x"963883ff",
   928 => x"f1b85275",
   929 => x"51811656",
   930 => x"8480808d",
   931 => x"a02d83ff",
   932 => x"f1b85780",
   933 => x"77848080",
   934 => x"80f52d56",
   935 => x"5474742e",
   936 => x"83388154",
   937 => x"7481e52e",
   938 => x"819c3881",
   939 => x"70750655",
   940 => x"5d73802e",
   941 => x"8190388b",
   942 => x"17848080",
   943 => x"80f52d98",
   944 => x"065b7a81",
   945 => x"81388b53",
   946 => x"7d527651",
   947 => x"84808092",
   948 => x"892d83ff",
   949 => x"e0800880",
   950 => x"ed389c17",
   951 => x"08518480",
   952 => x"808edd2d",
   953 => x"83ffe080",
   954 => x"08841d0c",
   955 => x"9a178480",
   956 => x"8080e02d",
   957 => x"51848080",
   958 => x"8f8f2d83",
   959 => x"ffe08008",
   960 => x"83ffe080",
   961 => x"08881e0c",
   962 => x"83ffe080",
   963 => x"08555583",
   964 => x"fff5dc08",
   965 => x"802ea038",
   966 => x"94178480",
   967 => x"8080e02d",
   968 => x"51848080",
   969 => x"8f8f2d83",
   970 => x"ffe08008",
   971 => x"902b83ff",
   972 => x"f00a0670",
   973 => x"16515473",
   974 => x"881d0c7a",
   975 => x"7c0c7c54",
   976 => x"8480809f",
   977 => x"a104811a",
   978 => x"5a848080",
   979 => x"9cee0483",
   980 => x"fff5dc08",
   981 => x"802e80c7",
   982 => x"38775184",
   983 => x"80809b8f",
   984 => x"2d83ffe0",
   985 => x"800883ff",
   986 => x"e0800853",
   987 => x"848080a6",
   988 => x"b8525884",
   989 => x"808082e3",
   990 => x"2d7780ff",
   991 => x"fffff806",
   992 => x"547380ff",
   993 => x"fffff82e",
   994 => x"9638fe18",
   995 => x"83fff5e4",
   996 => x"082983ff",
   997 => x"f5ec0805",
   998 => x"56848080",
   999 => x"9cec0480",
  1000 => x"547383ff",
  1001 => x"e0800c02",
  1002 => x"b8050d04",
  1003 => x"02f4050d",
  1004 => x"74700881",
  1005 => x"05710c70",
  1006 => x"0883fff5",
  1007 => x"d8080653",
  1008 => x"53719338",
  1009 => x"88130851",
  1010 => x"8480809b",
  1011 => x"8f2d83ff",
  1012 => x"e0800888",
  1013 => x"140c810b",
  1014 => x"83ffe080",
  1015 => x"0c028c05",
  1016 => x"0d0402f0",
  1017 => x"050d7588",
  1018 => x"1108fe05",
  1019 => x"83fff5e4",
  1020 => x"082983ff",
  1021 => x"f5ec0811",
  1022 => x"720883ff",
  1023 => x"f5d80806",
  1024 => x"05795553",
  1025 => x"54548480",
  1026 => x"808da02d",
  1027 => x"83ffe080",
  1028 => x"085383ff",
  1029 => x"e0800880",
  1030 => x"2e833881",
  1031 => x"537283ff",
  1032 => x"e0800c02",
  1033 => x"90050d04",
  1034 => x"02ec050d",
  1035 => x"76787154",
  1036 => x"83fff5bc",
  1037 => x"53545584",
  1038 => x"80809cb6",
  1039 => x"2d83ffe0",
  1040 => x"80085483",
  1041 => x"ffe08008",
  1042 => x"802e80ce",
  1043 => x"38848080",
  1044 => x"a6d05184",
  1045 => x"808085c5",
  1046 => x"2d83fff5",
  1047 => x"c00883ff",
  1048 => x"05892a55",
  1049 => x"80547375",
  1050 => x"2580d138",
  1051 => x"725283ff",
  1052 => x"f5bc5184",
  1053 => x"80809fe2",
  1054 => x"2d83ffe0",
  1055 => x"8008802e",
  1056 => x"af3883ff",
  1057 => x"f5bc5184",
  1058 => x"80809fac",
  1059 => x"2d848013",
  1060 => x"81155553",
  1061 => x"848080a0",
  1062 => x"e6047452",
  1063 => x"848080a6",
  1064 => x"ec518480",
  1065 => x"8082e32d",
  1066 => x"73538480",
  1067 => x"80a1be04",
  1068 => x"83ffe080",
  1069 => x"08538480",
  1070 => x"80a1be04",
  1071 => x"81537283",
  1072 => x"ffe0800c",
  1073 => x"0294050d",
  1074 => x"04000000",
  1075 => x"00ffffff",
  1076 => x"ff00ffff",
  1077 => x"ffff00ff",
  1078 => x"ffffff00",
  1079 => x"436d645f",
  1080 => x"696e6974",
  1081 => x"0a000000",
  1082 => x"636d645f",
  1083 => x"434d4438",
  1084 => x"20726573",
  1085 => x"706f6e73",
  1086 => x"653a2025",
  1087 => x"640a0000",
  1088 => x"434d4438",
  1089 => x"5f342072",
  1090 => x"6573706f",
  1091 => x"6e73653a",
  1092 => x"2025640a",
  1093 => x"00000000",
  1094 => x"53444843",
  1095 => x"20496e69",
  1096 => x"7469616c",
  1097 => x"697a6174",
  1098 => x"696f6e20",
  1099 => x"6572726f",
  1100 => x"72210a00",
  1101 => x"434d4435",
  1102 => x"38202564",
  1103 => x"0a202000",
  1104 => x"434d4435",
  1105 => x"385f3220",
  1106 => x"25640a20",
  1107 => x"20000000",
  1108 => x"53504920",
  1109 => x"496e6974",
  1110 => x"28290a00",
  1111 => x"52656164",
  1112 => x"20636f6d",
  1113 => x"6d616e64",
  1114 => x"20666169",
  1115 => x"6c656420",
  1116 => x"61742025",
  1117 => x"64202825",
  1118 => x"64290a00",
  1119 => x"496e6974",
  1120 => x"69616c69",
  1121 => x"7a696e67",
  1122 => x"20534420",
  1123 => x"63617264",
  1124 => x"0a000000",
  1125 => x"48756e74",
  1126 => x"696e6720",
  1127 => x"666f7220",
  1128 => x"70617274",
  1129 => x"6974696f",
  1130 => x"6e0a0000",
  1131 => x"4d414e49",
  1132 => x"46455354",
  1133 => x"4d535400",
  1134 => x"50617273",
  1135 => x"696e6720",
  1136 => x"6d616e69",
  1137 => x"66657374",
  1138 => x"0a000000",
  1139 => x"4c6f6164",
  1140 => x"696e6720",
  1141 => x"6d616e69",
  1142 => x"66657374",
  1143 => x"20666169",
  1144 => x"6c65640a",
  1145 => x"00000000",
  1146 => x"52657475",
  1147 => x"726e696e",
  1148 => x"670a0000",
  1149 => x"52656164",
  1150 => x"696e6720",
  1151 => x"4d42520a",
  1152 => x"00000000",
  1153 => x"52656164",
  1154 => x"206f6620",
  1155 => x"4d425220",
  1156 => x"6661696c",
  1157 => x"65640a00",
  1158 => x"4d425220",
  1159 => x"73756363",
  1160 => x"65737366",
  1161 => x"756c6c79",
  1162 => x"20726561",
  1163 => x"640a0000",
  1164 => x"46415431",
  1165 => x"36202020",
  1166 => x"00000000",
  1167 => x"46415433",
  1168 => x"32202020",
  1169 => x"00000000",
  1170 => x"50617274",
  1171 => x"6974696f",
  1172 => x"6e636f75",
  1173 => x"6e742025",
  1174 => x"640a0000",
  1175 => x"4e6f2070",
  1176 => x"61727469",
  1177 => x"74696f6e",
  1178 => x"20736967",
  1179 => x"6e617475",
  1180 => x"72652066",
  1181 => x"6f756e64",
  1182 => x"0a000000",
  1183 => x"52656164",
  1184 => x"696e6720",
  1185 => x"626f6f74",
  1186 => x"20736563",
  1187 => x"746f7220",
  1188 => x"25640a00",
  1189 => x"52656164",
  1190 => x"20626f6f",
  1191 => x"74207365",
  1192 => x"63746f72",
  1193 => x"2066726f",
  1194 => x"6d206669",
  1195 => x"72737420",
  1196 => x"70617274",
  1197 => x"6974696f",
  1198 => x"6e0a0000",
  1199 => x"48756e74",
  1200 => x"696e6720",
  1201 => x"666f7220",
  1202 => x"66696c65",
  1203 => x"73797374",
  1204 => x"656d0a00",
  1205 => x"556e7375",
  1206 => x"70706f72",
  1207 => x"74656420",
  1208 => x"70617274",
  1209 => x"6974696f",
  1210 => x"6e207479",
  1211 => x"7065210d",
  1212 => x"00000000",
  1213 => x"436c7573",
  1214 => x"74657220",
  1215 => x"73697a65",
  1216 => x"3a202564",
  1217 => x"2c20436c",
  1218 => x"75737465",
  1219 => x"72206d61",
  1220 => x"736b2c20",
  1221 => x"25640a00",
  1222 => x"47657443",
  1223 => x"6c757374",
  1224 => x"65722072",
  1225 => x"65616469",
  1226 => x"6e672073",
  1227 => x"6563746f",
  1228 => x"72202564",
  1229 => x"0a000000",
  1230 => x"47657446",
  1231 => x"41544c69",
  1232 => x"6e6b2072",
  1233 => x"65747572",
  1234 => x"6e656420",
  1235 => x"25640a00",
  1236 => x"4f70656e",
  1237 => x"65642066",
  1238 => x"696c652c",
  1239 => x"206c6f61",
  1240 => x"64696e67",
  1241 => x"2e2e2e0a",
  1242 => x"00000000",
  1243 => x"43616e27",
  1244 => x"74206f70",
  1245 => x"656e2025",
  1246 => x"730a0000",
	others => x"00000000"
);

begin

process (clk)
begin
	if (clk'event and clk = '1') then
		if (from_zpu.memAWriteEnable = '1') and (from_zpu.memBWriteEnable = '1') and (from_zpu.memAAddr=from_zpu.memBAddr) and (from_zpu.memAWrite/=from_zpu.memBWrite) then
			report "write collision" severity failure;
		end if;
	
		if (from_zpu.memAWriteEnable = '1') then
			ram(to_integer(unsigned(from_zpu.memAAddr(maxAddrBitBRAM downto 2)))) := from_zpu.memAWrite;
			to_zpu.memARead <= from_zpu.memAWrite;
		else
			to_zpu.memARead <= ram(to_integer(unsigned(from_zpu.memAAddr(maxAddrBitBRAM downto 2))));
		end if;
	end if;
end process;

process (clk)
begin
	if (clk'event and clk = '1') then
		if (from_zpu.memBWriteEnable = '1') then
			ram(to_integer(unsigned(from_zpu.memBAddr(maxAddrBitBRAM downto 2)))) := from_zpu.memBWrite;
			to_zpu.memBRead <= from_zpu.memBWrite;
		else
			to_zpu.memBRead <= ram(to_integer(unsigned(from_zpu.memBAddr(maxAddrBitBRAM downto 2))));
		end if;
	end if;
end process;


end arch;

