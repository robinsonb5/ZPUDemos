-- ZPU
--
-- Copyright 2004-2008 oharboe - �yvind Harboe - oyvind.harboe@zylin.com
-- Modified by Alastair M. Robinson for the ZPUFlex project.
--
-- The FreeBSD license
-- 
-- Redistribution and use in source and binary forms, with or without
-- modification, are permitted provided that the following conditions
-- are met:
-- 
-- 1. Redistributions of source code must retain the above copyright
--    notice, this list of conditions and the following disclaimer.
-- 2. Redistributions in binary form must reproduce the above
--    copyright notice, this list of conditions and the following
--    disclaimer in the documentation and/or other materials
--    provided with the distribution.
-- 
-- THIS SOFTWARE IS PROVIDED BY THE ZPU PROJECT ``AS IS'' AND ANY
-- EXPRESS OR IMPLIED WARRANTIES, INCLUDING, BUT NOT LIMITED TO,
-- THE IMPLIED WARRANTIES OF MERCHANTABILITY AND FITNESS FOR A
-- PARTICULAR PURPOSE ARE DISCLAIMED. IN NO EVENT SHALL THE
-- ZPU PROJECT OR CONTRIBUTORS BE LIABLE FOR ANY DIRECT,
-- INDIRECT, INCIDENTAL, SPECIAL, EXEMPLARY, OR CONSEQUENTIAL DAMAGES
-- (INCLUDING, BUT NOT LIMITED TO, PROCUREMENT OF SUBSTITUTE GOODS
-- OR SERVICES; LOSS OF USE, DATA, OR PROFITS; OR BUSINESS INTERRUPTION)
-- HOWEVER CAUSED AND ON ANY THEORY OF LIABILITY, WHETHER IN CONTRACT,
-- STRICT LIABILITY, OR TORT (INCLUDING NEGLIGENCE OR OTHERWISE)
-- ARISING IN ANY WAY OUT OF THE USE OF THIS SOFTWARE, EVEN IF
-- ADVISED OF THE POSSIBILITY OF SUCH DAMAGE.
-- 
-- The views and conclusions contained in the software and documentation
-- are those of the authors and should not be interpreted as representing
-- official policies, either expressed or implied, of the ZPU Project.

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;


library work;
use work.zpu_config.all;
use work.zpupkg.all;

entity Dhrystone_min_ROM is
generic
	(
		maxAddrBit : integer := maxAddrBitBRAMLimit -- Specify your actual ROM size to save LEs and unnecessary block RAM usage.
	);
port (
	clk : in std_logic;
	areset : in std_logic := '0';
	from_zpu : in ZPU_ToROM;
	to_zpu : out ZPU_FromROM
);
end Dhrystone_min_ROM;

architecture arch of Dhrystone_min_ROM is

type ram_type is array(natural range 0 to ((2**(maxAddrBit+1))/4)-1) of std_logic_vector(wordSize-1 downto 0);

shared variable ram : ram_type :=
(
     0 => x"0b0b0b88",
     1 => x"dd040000",
     2 => x"00000000",
     3 => x"00000000",
     4 => x"00000000",
     5 => x"00000000",
     6 => x"00000000",
     7 => x"00000000",
     8 => x"04000000",
     9 => x"00000000",
    10 => x"00000000",
    11 => x"00000000",
    12 => x"00000000",
    13 => x"00000000",
    14 => x"00000000",
    15 => x"00000000",
    16 => x"71fd0608",
    17 => x"72830609",
    18 => x"81058205",
    19 => x"832b2a83",
    20 => x"ffff0652",
    21 => x"04000000",
    22 => x"00000000",
    23 => x"00000000",
    24 => x"71fd0608",
    25 => x"83ffff73",
    26 => x"83060981",
    27 => x"05820583",
    28 => x"2b2b0906",
    29 => x"7383ffff",
    30 => x"0b0b0b0b",
    31 => x"83a50400",
    32 => x"72098105",
    33 => x"72057373",
    34 => x"09060906",
    35 => x"73097306",
    36 => x"070a8106",
    37 => x"53510400",
    38 => x"00000000",
    39 => x"00000000",
    40 => x"72722473",
    41 => x"732e0753",
    42 => x"51040000",
    43 => x"00000000",
    44 => x"00000000",
    45 => x"00000000",
    46 => x"00000000",
    47 => x"00000000",
    48 => x"71737109",
    49 => x"71068106",
    50 => x"09810572",
    51 => x"0a100a72",
    52 => x"0a100a31",
    53 => x"050a8106",
    54 => x"51515351",
    55 => x"04000000",
    56 => x"72722673",
    57 => x"732e0753",
    58 => x"51040000",
    59 => x"00000000",
    60 => x"00000000",
    61 => x"00000000",
    62 => x"00000000",
    63 => x"00000000",
    64 => x"00000000",
    65 => x"00000000",
    66 => x"00000000",
    67 => x"00000000",
    68 => x"00000000",
    69 => x"00000000",
    70 => x"00000000",
    71 => x"00000000",
    72 => x"0b0b0b88",
    73 => x"ba040000",
    74 => x"00000000",
    75 => x"00000000",
    76 => x"00000000",
    77 => x"00000000",
    78 => x"00000000",
    79 => x"00000000",
    80 => x"720a722b",
    81 => x"0a535104",
    82 => x"00000000",
    83 => x"00000000",
    84 => x"00000000",
    85 => x"00000000",
    86 => x"00000000",
    87 => x"00000000",
    88 => x"72729f06",
    89 => x"0981050b",
    90 => x"0b0b889f",
    91 => x"05040000",
    92 => x"00000000",
    93 => x"00000000",
    94 => x"00000000",
    95 => x"00000000",
    96 => x"72722aff",
    97 => x"739f062a",
    98 => x"0974090a",
    99 => x"8106ff05",
   100 => x"06075351",
   101 => x"04000000",
   102 => x"00000000",
   103 => x"00000000",
   104 => x"71715351",
   105 => x"04067383",
   106 => x"06098105",
   107 => x"8205832b",
   108 => x"0b2b0772",
   109 => x"fc060c51",
   110 => x"51040000",
   111 => x"00000000",
   112 => x"72098105",
   113 => x"72050970",
   114 => x"81050906",
   115 => x"0a810653",
   116 => x"51040000",
   117 => x"00000000",
   118 => x"00000000",
   119 => x"00000000",
   120 => x"72098105",
   121 => x"72050970",
   122 => x"81050906",
   123 => x"0a098106",
   124 => x"53510400",
   125 => x"00000000",
   126 => x"00000000",
   127 => x"00000000",
   128 => x"71098105",
   129 => x"52040000",
   130 => x"00000000",
   131 => x"00000000",
   132 => x"00000000",
   133 => x"00000000",
   134 => x"00000000",
   135 => x"00000000",
   136 => x"72720981",
   137 => x"05055351",
   138 => x"04000000",
   139 => x"00000000",
   140 => x"00000000",
   141 => x"00000000",
   142 => x"00000000",
   143 => x"00000000",
   144 => x"72097206",
   145 => x"73730906",
   146 => x"07535104",
   147 => x"00000000",
   148 => x"00000000",
   149 => x"00000000",
   150 => x"00000000",
   151 => x"00000000",
   152 => x"71fc0608",
   153 => x"72830609",
   154 => x"81058305",
   155 => x"1010102a",
   156 => x"81ff0652",
   157 => x"04000000",
   158 => x"00000000",
   159 => x"00000000",
   160 => x"71fc0608",
   161 => x"0b0b0b9f",
   162 => x"e8738306",
   163 => x"10100508",
   164 => x"060b0b0b",
   165 => x"88a20400",
   166 => x"00000000",
   167 => x"00000000",
   168 => x"88088c08",
   169 => x"90087575",
   170 => x"0b0b0b98",
   171 => x"db2d5050",
   172 => x"88085690",
   173 => x"0c8c0c88",
   174 => x"0c510400",
   175 => x"00000000",
   176 => x"88088c08",
   177 => x"90087575",
   178 => x"0b0b0b9a",
   179 => x"8d2d5050",
   180 => x"88085690",
   181 => x"0c8c0c88",
   182 => x"0c510400",
   183 => x"00000000",
   184 => x"72097081",
   185 => x"0509060a",
   186 => x"8106ff05",
   187 => x"70547106",
   188 => x"73097274",
   189 => x"05ff0506",
   190 => x"07515151",
   191 => x"04000000",
   192 => x"72097081",
   193 => x"0509060a",
   194 => x"098106ff",
   195 => x"05705471",
   196 => x"06730972",
   197 => x"7405ff05",
   198 => x"06075151",
   199 => x"51040000",
   200 => x"05ff0504",
   201 => x"00000000",
   202 => x"00000000",
   203 => x"00000000",
   204 => x"00000000",
   205 => x"00000000",
   206 => x"00000000",
   207 => x"00000000",
   208 => x"04000000",
   209 => x"00000000",
   210 => x"00000000",
   211 => x"00000000",
   212 => x"00000000",
   213 => x"00000000",
   214 => x"00000000",
   215 => x"00000000",
   216 => x"71810552",
   217 => x"04000000",
   218 => x"00000000",
   219 => x"00000000",
   220 => x"00000000",
   221 => x"00000000",
   222 => x"00000000",
   223 => x"00000000",
   224 => x"00000000",
   225 => x"00000000",
   226 => x"00000000",
   227 => x"00000000",
   228 => x"00000000",
   229 => x"00000000",
   230 => x"00000000",
   231 => x"00000000",
   232 => x"02840572",
   233 => x"10100552",
   234 => x"04000000",
   235 => x"00000000",
   236 => x"00000000",
   237 => x"00000000",
   238 => x"00000000",
   239 => x"00000000",
   240 => x"00000000",
   241 => x"00000000",
   242 => x"00000000",
   243 => x"00000000",
   244 => x"00000000",
   245 => x"00000000",
   246 => x"00000000",
   247 => x"00000000",
   248 => x"717105ff",
   249 => x"05715351",
   250 => x"020d0400",
   251 => x"00000000",
   252 => x"00000000",
   253 => x"00000000",
   254 => x"00000000",
   255 => x"00000000",
   256 => x"10101010",
   257 => x"10101010",
   258 => x"10101010",
   259 => x"10101010",
   260 => x"10101010",
   261 => x"10101010",
   262 => x"10101010",
   263 => x"10101053",
   264 => x"51047381",
   265 => x"ff067383",
   266 => x"06098105",
   267 => x"83051010",
   268 => x"102b0772",
   269 => x"fc060c51",
   270 => x"51047272",
   271 => x"80728106",
   272 => x"ff050972",
   273 => x"06057110",
   274 => x"52720a10",
   275 => x"0a5372ed",
   276 => x"38515153",
   277 => x"51040000",
   278 => x"800488da",
   279 => x"0488da0b",
   280 => x"8ef004f1",
   281 => x"3d0d923d",
   282 => x"0b0b0ba5",
   283 => x"905a5c80",
   284 => x"7c708405",
   285 => x"5e08715f",
   286 => x"5f577d70",
   287 => x"84055f08",
   288 => x"56805875",
   289 => x"982a7688",
   290 => x"2b575574",
   291 => x"802e82b8",
   292 => x"387c802e",
   293 => x"b738805d",
   294 => x"7480e42e",
   295 => x"81983874",
   296 => x"80e42680",
   297 => x"d8387480",
   298 => x"e32eb738",
   299 => x"a551829f",
   300 => x"3f745182",
   301 => x"9a3f8217",
   302 => x"57811858",
   303 => x"837825c3",
   304 => x"3874ffb6",
   305 => x"387e880c",
   306 => x"913d0d04",
   307 => x"74a52e09",
   308 => x"81069738",
   309 => x"810b8119",
   310 => x"595d8378",
   311 => x"25ffa438",
   312 => x"e0397b84",
   313 => x"1d710857",
   314 => x"5d5a7451",
   315 => x"81e13f81",
   316 => x"17811959",
   317 => x"57837825",
   318 => x"ff8938c5",
   319 => x"397480f3",
   320 => x"2e098106",
   321 => x"ffa6387b",
   322 => x"841d7108",
   323 => x"70545b5d",
   324 => x"5481db3f",
   325 => x"800bff11",
   326 => x"55538073",
   327 => x"25ff9a38",
   328 => x"78708105",
   329 => x"5a337052",
   330 => x"5581a43f",
   331 => x"811774ff",
   332 => x"16565457",
   333 => x"e5397b84",
   334 => x"1d71080b",
   335 => x"0b0ba590",
   336 => x"0b0b0b0b",
   337 => x"a4c0615f",
   338 => x"585e525d",
   339 => x"5372b138",
   340 => x"b00b0b0b",
   341 => x"0ba4c034",
   342 => x"811454ff",
   343 => x"14547333",
   344 => x"7b708105",
   345 => x"5d34811a",
   346 => x"5a730b0b",
   347 => x"0ba4c02e",
   348 => x"098106e7",
   349 => x"38807b34",
   350 => x"79ff1155",
   351 => x"53ff9b39",
   352 => x"8a527251",
   353 => x"8db03f88",
   354 => x"080b0b0b",
   355 => x"9ff80533",
   356 => x"74708105",
   357 => x"56348a52",
   358 => x"72518cf5",
   359 => x"3f880853",
   360 => x"8808dd38",
   361 => x"730b0b0b",
   362 => x"a4c02ec9",
   363 => x"38ff1454",
   364 => x"73337b70",
   365 => x"81055d34",
   366 => x"811a5a73",
   367 => x"0b0b0ba4",
   368 => x"c02effb1",
   369 => x"38ff9439",
   370 => x"76880c91",
   371 => x"3d0d04ff",
   372 => x"3d0d7352",
   373 => x"c0087088",
   374 => x"2a708106",
   375 => x"51515170",
   376 => x"802ef138",
   377 => x"71c00c71",
   378 => x"880c833d",
   379 => x"0d04fb3d",
   380 => x"0d775675",
   381 => x"70840557",
   382 => x"08538054",
   383 => x"72982a73",
   384 => x"882b5452",
   385 => x"71802ea2",
   386 => x"38c00870",
   387 => x"882a7081",
   388 => x"06515151",
   389 => x"70802ef1",
   390 => x"3871c00c",
   391 => x"81158115",
   392 => x"55558374",
   393 => x"25d63871",
   394 => x"ca387488",
   395 => x"0c873d0d",
   396 => x"04c80888",
   397 => x"0c04803d",
   398 => x"0d80c10b",
   399 => x"80f4dc34",
   400 => x"800b80f6",
   401 => x"f40c7088",
   402 => x"0c823d0d",
   403 => x"04ff3d0d",
   404 => x"800b80f4",
   405 => x"dc335252",
   406 => x"7080c12e",
   407 => x"99387180",
   408 => x"f6f40807",
   409 => x"80f6f40c",
   410 => x"80c20b80",
   411 => x"f4e03470",
   412 => x"880c833d",
   413 => x"0d04810b",
   414 => x"80f6f408",
   415 => x"0780f6f4",
   416 => x"0c80c20b",
   417 => x"80f4e034",
   418 => x"70880c83",
   419 => x"3d0d04fd",
   420 => x"3d0d7570",
   421 => x"088a0553",
   422 => x"5380f4dc",
   423 => x"33517080",
   424 => x"c12e8b38",
   425 => x"73f33870",
   426 => x"880c853d",
   427 => x"0d04ff12",
   428 => x"7080f4d8",
   429 => x"0831740c",
   430 => x"880c853d",
   431 => x"0d04fc3d",
   432 => x"0d80f584",
   433 => x"08557480",
   434 => x"2e8c3876",
   435 => x"7508710c",
   436 => x"80f58408",
   437 => x"56548c15",
   438 => x"5380f4d8",
   439 => x"08528a51",
   440 => x"889c3f73",
   441 => x"880c863d",
   442 => x"0d04fb3d",
   443 => x"0d777008",
   444 => x"5656b053",
   445 => x"80f58408",
   446 => x"5274518f",
   447 => x"bc3f850b",
   448 => x"8c170c85",
   449 => x"0b8c160c",
   450 => x"7508750c",
   451 => x"80f58408",
   452 => x"5473802e",
   453 => x"8a387308",
   454 => x"750c80f5",
   455 => x"8408548c",
   456 => x"145380f4",
   457 => x"d808528a",
   458 => x"5187d33f",
   459 => x"841508ad",
   460 => x"38860b8c",
   461 => x"160c8815",
   462 => x"52881608",
   463 => x"5186df3f",
   464 => x"80f58408",
   465 => x"7008760c",
   466 => x"548c1570",
   467 => x"54548a52",
   468 => x"73085187",
   469 => x"a93f7388",
   470 => x"0c873d0d",
   471 => x"04750854",
   472 => x"b0537352",
   473 => x"75518ed1",
   474 => x"3f73880c",
   475 => x"873d0d04",
   476 => x"f33d0d80",
   477 => x"f3f00b80",
   478 => x"f4a40c80",
   479 => x"f4a80b80",
   480 => x"f5840c80",
   481 => x"f3f00b80",
   482 => x"f4a80c80",
   483 => x"0b80f4a8",
   484 => x"0b84050c",
   485 => x"820b80f4",
   486 => x"a80b8805",
   487 => x"0ca80b80",
   488 => x"f4a80b8c",
   489 => x"050c9f53",
   490 => x"a08c5280",
   491 => x"f4b8518e",
   492 => x"883f9f53",
   493 => x"a0ac5280",
   494 => x"f6d4518d",
   495 => x"fc3f8a0b",
   496 => x"b2bc0ca3",
   497 => x"8c51f99b",
   498 => x"3fa0cc51",
   499 => x"f9953fa3",
   500 => x"8c51f98f",
   501 => x"3fa4bc08",
   502 => x"802e83e6",
   503 => x"38a0fc51",
   504 => x"f9813fa3",
   505 => x"8c51f8fb",
   506 => x"3fa4b808",
   507 => x"52a1a851",
   508 => x"f8f13fc8",
   509 => x"0870a5dc",
   510 => x"0c568158",
   511 => x"800ba4b8",
   512 => x"082582c4",
   513 => x"388c3d5b",
   514 => x"80c10b80",
   515 => x"f4dc3481",
   516 => x"0b80f6f4",
   517 => x"0c80c20b",
   518 => x"80f4e034",
   519 => x"825c835a",
   520 => x"9f53a1d8",
   521 => x"5280f4e4",
   522 => x"518d8e3f",
   523 => x"815d800b",
   524 => x"80f4e453",
   525 => x"80f6d452",
   526 => x"5586e73f",
   527 => x"8808752e",
   528 => x"09810683",
   529 => x"38815574",
   530 => x"80f6f40c",
   531 => x"7b705755",
   532 => x"748325a0",
   533 => x"38741010",
   534 => x"15fd055e",
   535 => x"8f3dfc05",
   536 => x"53835275",
   537 => x"5185973f",
   538 => x"811c705d",
   539 => x"70575583",
   540 => x"7524e238",
   541 => x"7d547453",
   542 => x"a5e05280",
   543 => x"f58c5185",
   544 => x"8d3f80f5",
   545 => x"84087008",
   546 => x"5757b053",
   547 => x"76527551",
   548 => x"8ca73f85",
   549 => x"0b8c180c",
   550 => x"850b8c17",
   551 => x"0c760876",
   552 => x"0c80f584",
   553 => x"08557480",
   554 => x"2e8a3874",
   555 => x"08760c80",
   556 => x"f5840855",
   557 => x"8c155380",
   558 => x"f4d80852",
   559 => x"8a5184be",
   560 => x"3f841608",
   561 => x"839e3886",
   562 => x"0b8c170c",
   563 => x"88165288",
   564 => x"17085183",
   565 => x"c93f80f5",
   566 => x"84087008",
   567 => x"770c578c",
   568 => x"16705455",
   569 => x"8a527408",
   570 => x"5184933f",
   571 => x"80c10b80",
   572 => x"f4e03356",
   573 => x"56757526",
   574 => x"a23880c3",
   575 => x"52755184",
   576 => x"f73f8808",
   577 => x"7d2e82af",
   578 => x"38811670",
   579 => x"81ff0680",
   580 => x"f4e03352",
   581 => x"57557476",
   582 => x"27e0387d",
   583 => x"7a7d2935",
   584 => x"705d8a05",
   585 => x"80f4dc33",
   586 => x"80f4d808",
   587 => x"59575575",
   588 => x"80c12e82",
   589 => x"c73878f7",
   590 => x"38811858",
   591 => x"a4b80878",
   592 => x"25fdc538",
   593 => x"a5dc0856",
   594 => x"c8087080",
   595 => x"f4a00c70",
   596 => x"773170a5",
   597 => x"d80c53a1",
   598 => x"f8525bf6",
   599 => x"863fa5d8",
   600 => x"085680f7",
   601 => x"762580e0",
   602 => x"38a4b808",
   603 => x"707787e8",
   604 => x"2935a5d0",
   605 => x"0c767187",
   606 => x"e82935a5",
   607 => x"d40c7671",
   608 => x"84b92935",
   609 => x"80f5880c",
   610 => x"5aa28851",
   611 => x"f5d53fa5",
   612 => x"d00852a2",
   613 => x"b851f5cb",
   614 => x"3fa2c051",
   615 => x"f5c53fa5",
   616 => x"d40852a2",
   617 => x"b851f5bb",
   618 => x"3f80f588",
   619 => x"0852a2f0",
   620 => x"51f5b03f",
   621 => x"a38c51f5",
   622 => x"aa3f800b",
   623 => x"880c8f3d",
   624 => x"0d04a390",
   625 => x"51fc9939",
   626 => x"a3c051f5",
   627 => x"963fa3f8",
   628 => x"51f5903f",
   629 => x"a38c51f5",
   630 => x"8a3fa5d8",
   631 => x"08a4b808",
   632 => x"707287e8",
   633 => x"2935a5d0",
   634 => x"0c717187",
   635 => x"e82935a5",
   636 => x"d40c7171",
   637 => x"84b92935",
   638 => x"80f5880c",
   639 => x"5b56a288",
   640 => x"51f4e03f",
   641 => x"a5d00852",
   642 => x"a2b851f4",
   643 => x"d63fa2c0",
   644 => x"51f4d03f",
   645 => x"a5d40852",
   646 => x"a2b851f4",
   647 => x"c63f80f5",
   648 => x"880852a2",
   649 => x"f051f4bb",
   650 => x"3fa38c51",
   651 => x"f4b53f80",
   652 => x"0b880c8f",
   653 => x"3d0d048f",
   654 => x"3df80552",
   655 => x"805180de",
   656 => x"3f9f53a4",
   657 => x"985280f4",
   658 => x"e45188ed",
   659 => x"3f777880",
   660 => x"f4d80c81",
   661 => x"177081ff",
   662 => x"0680f4e0",
   663 => x"33525856",
   664 => x"5afdb339",
   665 => x"760856b0",
   666 => x"53755276",
   667 => x"5188ca3f",
   668 => x"80c10b80",
   669 => x"f4e03356",
   670 => x"56fcfa39",
   671 => x"ff157078",
   672 => x"317c0c59",
   673 => x"8059fdb1",
   674 => x"39ff3d0d",
   675 => x"73823270",
   676 => x"30707207",
   677 => x"8025880c",
   678 => x"5252833d",
   679 => x"0d04fe3d",
   680 => x"0d747671",
   681 => x"53545271",
   682 => x"822e8338",
   683 => x"83517181",
   684 => x"2e9a3881",
   685 => x"72269f38",
   686 => x"71822eb8",
   687 => x"3871842e",
   688 => x"a9387073",
   689 => x"0c70880c",
   690 => x"843d0d04",
   691 => x"80e40b80",
   692 => x"f4d80825",
   693 => x"8b388073",
   694 => x"0c70880c",
   695 => x"843d0d04",
   696 => x"83730c70",
   697 => x"880c843d",
   698 => x"0d048273",
   699 => x"0c70880c",
   700 => x"843d0d04",
   701 => x"81730c70",
   702 => x"880c843d",
   703 => x"0d04803d",
   704 => x"0d747414",
   705 => x"8205710c",
   706 => x"880c823d",
   707 => x"0d04f73d",
   708 => x"0d7b7d7f",
   709 => x"61851270",
   710 => x"822b7511",
   711 => x"70747170",
   712 => x"8405530c",
   713 => x"5a5a5d5b",
   714 => x"760c7980",
   715 => x"f8180c79",
   716 => x"86125257",
   717 => x"585a5a76",
   718 => x"76249938",
   719 => x"76b32982",
   720 => x"2b791151",
   721 => x"53767370",
   722 => x"8405550c",
   723 => x"81145475",
   724 => x"7425f238",
   725 => x"7681cc29",
   726 => x"19fc1108",
   727 => x"8105fc12",
   728 => x"0c7a1970",
   729 => x"089fa013",
   730 => x"0c585685",
   731 => x"0b80f4d8",
   732 => x"0c75880c",
   733 => x"8b3d0d04",
   734 => x"fe3d0d02",
   735 => x"93053351",
   736 => x"80028405",
   737 => x"97053354",
   738 => x"5270732e",
   739 => x"88387188",
   740 => x"0c843d0d",
   741 => x"047080f4",
   742 => x"dc34810b",
   743 => x"880c843d",
   744 => x"0d04f83d",
   745 => x"0d7a7c59",
   746 => x"56820b83",
   747 => x"19555574",
   748 => x"16703375",
   749 => x"335b5153",
   750 => x"72792e80",
   751 => x"c63880c1",
   752 => x"0b811681",
   753 => x"16565657",
   754 => x"827525e3",
   755 => x"38ffa917",
   756 => x"7081ff06",
   757 => x"55597382",
   758 => x"26833887",
   759 => x"55815376",
   760 => x"80d22e98",
   761 => x"38775275",
   762 => x"5186e73f",
   763 => x"80537288",
   764 => x"08258938",
   765 => x"871580f4",
   766 => x"d80c8153",
   767 => x"72880c8a",
   768 => x"3d0d0472",
   769 => x"80f4dc34",
   770 => x"827525ff",
   771 => x"a238ffbd",
   772 => x"39940802",
   773 => x"940cfd3d",
   774 => x"0d805394",
   775 => x"088c0508",
   776 => x"52940888",
   777 => x"05085182",
   778 => x"de3f8808",
   779 => x"70880c54",
   780 => x"853d0d94",
   781 => x"0c049408",
   782 => x"02940cfd",
   783 => x"3d0d8153",
   784 => x"94088c05",
   785 => x"08529408",
   786 => x"88050851",
   787 => x"82b93f88",
   788 => x"0870880c",
   789 => x"54853d0d",
   790 => x"940c0494",
   791 => x"0802940c",
   792 => x"f93d0d80",
   793 => x"0b9408fc",
   794 => x"050c9408",
   795 => x"88050880",
   796 => x"25ab3894",
   797 => x"08880508",
   798 => x"30940888",
   799 => x"050c800b",
   800 => x"9408f405",
   801 => x"0c9408fc",
   802 => x"05088838",
   803 => x"810b9408",
   804 => x"f4050c94",
   805 => x"08f40508",
   806 => x"9408fc05",
   807 => x"0c94088c",
   808 => x"05088025",
   809 => x"ab389408",
   810 => x"8c050830",
   811 => x"94088c05",
   812 => x"0c800b94",
   813 => x"08f0050c",
   814 => x"9408fc05",
   815 => x"08883881",
   816 => x"0b9408f0",
   817 => x"050c9408",
   818 => x"f0050894",
   819 => x"08fc050c",
   820 => x"80539408",
   821 => x"8c050852",
   822 => x"94088805",
   823 => x"085181a7",
   824 => x"3f880870",
   825 => x"9408f805",
   826 => x"0c549408",
   827 => x"fc050880",
   828 => x"2e8c3894",
   829 => x"08f80508",
   830 => x"309408f8",
   831 => x"050c9408",
   832 => x"f8050870",
   833 => x"880c5489",
   834 => x"3d0d940c",
   835 => x"04940802",
   836 => x"940cfb3d",
   837 => x"0d800b94",
   838 => x"08fc050c",
   839 => x"94088805",
   840 => x"08802593",
   841 => x"38940888",
   842 => x"05083094",
   843 => x"0888050c",
   844 => x"810b9408",
   845 => x"fc050c94",
   846 => x"088c0508",
   847 => x"80258c38",
   848 => x"94088c05",
   849 => x"08309408",
   850 => x"8c050c81",
   851 => x"5394088c",
   852 => x"05085294",
   853 => x"08880508",
   854 => x"51ad3f88",
   855 => x"08709408",
   856 => x"f8050c54",
   857 => x"9408fc05",
   858 => x"08802e8c",
   859 => x"389408f8",
   860 => x"05083094",
   861 => x"08f8050c",
   862 => x"9408f805",
   863 => x"0870880c",
   864 => x"54873d0d",
   865 => x"940c0494",
   866 => x"0802940c",
   867 => x"fd3d0d81",
   868 => x"0b9408fc",
   869 => x"050c800b",
   870 => x"9408f805",
   871 => x"0c94088c",
   872 => x"05089408",
   873 => x"88050827",
   874 => x"ac389408",
   875 => x"fc050880",
   876 => x"2ea33880",
   877 => x"0b94088c",
   878 => x"05082499",
   879 => x"3894088c",
   880 => x"05081094",
   881 => x"088c050c",
   882 => x"9408fc05",
   883 => x"08109408",
   884 => x"fc050cc9",
   885 => x"399408fc",
   886 => x"0508802e",
   887 => x"80c93894",
   888 => x"088c0508",
   889 => x"94088805",
   890 => x"0826a138",
   891 => x"94088805",
   892 => x"0894088c",
   893 => x"05083194",
   894 => x"0888050c",
   895 => x"9408f805",
   896 => x"089408fc",
   897 => x"05080794",
   898 => x"08f8050c",
   899 => x"9408fc05",
   900 => x"08812a94",
   901 => x"08fc050c",
   902 => x"94088c05",
   903 => x"08812a94",
   904 => x"088c050c",
   905 => x"ffaf3994",
   906 => x"08900508",
   907 => x"802e8f38",
   908 => x"94088805",
   909 => x"08709408",
   910 => x"f4050c51",
   911 => x"8d399408",
   912 => x"f8050870",
   913 => x"9408f405",
   914 => x"0c519408",
   915 => x"f4050888",
   916 => x"0c853d0d",
   917 => x"940c0494",
   918 => x"0802940c",
   919 => x"ff3d0d80",
   920 => x"0b9408fc",
   921 => x"050c9408",
   922 => x"88050881",
   923 => x"06ff1170",
   924 => x"09709408",
   925 => x"8c050806",
   926 => x"9408fc05",
   927 => x"08119408",
   928 => x"fc050c94",
   929 => x"08880508",
   930 => x"812a9408",
   931 => x"88050c94",
   932 => x"088c0508",
   933 => x"1094088c",
   934 => x"050c5151",
   935 => x"51519408",
   936 => x"88050880",
   937 => x"2e8438ff",
   938 => x"bd399408",
   939 => x"fc050870",
   940 => x"880c5183",
   941 => x"3d0d940c",
   942 => x"04fc3d0d",
   943 => x"7670797b",
   944 => x"55555555",
   945 => x"8f72278c",
   946 => x"38727507",
   947 => x"83065170",
   948 => x"802ea738",
   949 => x"ff125271",
   950 => x"ff2e9838",
   951 => x"72708105",
   952 => x"54337470",
   953 => x"81055634",
   954 => x"ff125271",
   955 => x"ff2e0981",
   956 => x"06ea3874",
   957 => x"880c863d",
   958 => x"0d047451",
   959 => x"72708405",
   960 => x"54087170",
   961 => x"8405530c",
   962 => x"72708405",
   963 => x"54087170",
   964 => x"8405530c",
   965 => x"72708405",
   966 => x"54087170",
   967 => x"8405530c",
   968 => x"72708405",
   969 => x"54087170",
   970 => x"8405530c",
   971 => x"f0125271",
   972 => x"8f26c938",
   973 => x"83722795",
   974 => x"38727084",
   975 => x"05540871",
   976 => x"70840553",
   977 => x"0cfc1252",
   978 => x"718326ed",
   979 => x"387054ff",
   980 => x"8339fb3d",
   981 => x"0d777970",
   982 => x"72078306",
   983 => x"53545270",
   984 => x"93387173",
   985 => x"73085456",
   986 => x"54717308",
   987 => x"2e80c438",
   988 => x"73755452",
   989 => x"71337081",
   990 => x"ff065254",
   991 => x"70802e9d",
   992 => x"38723355",
   993 => x"70752e09",
   994 => x"81069538",
   995 => x"81128114",
   996 => x"71337081",
   997 => x"ff065456",
   998 => x"545270e5",
   999 => x"38723355",
  1000 => x"7381ff06",
  1001 => x"7581ff06",
  1002 => x"71713188",
  1003 => x"0c525287",
  1004 => x"3d0d0471",
  1005 => x"0970f7fb",
  1006 => x"fdff1406",
  1007 => x"70f88482",
  1008 => x"81800651",
  1009 => x"51517097",
  1010 => x"38841484",
  1011 => x"16710854",
  1012 => x"56547175",
  1013 => x"082edc38",
  1014 => x"73755452",
  1015 => x"ff963980",
  1016 => x"0b880c87",
  1017 => x"3d0d0400",
  1018 => x"00ffffff",
  1019 => x"ff00ffff",
  1020 => x"ffff00ff",
  1021 => x"ffffff00",
  1022 => x"30313233",
  1023 => x"34353637",
  1024 => x"38394142",
  1025 => x"43444546",
  1026 => x"00000000",
  1027 => x"44485259",
  1028 => x"53544f4e",
  1029 => x"45205052",
  1030 => x"4f475241",
  1031 => x"4d2c2053",
  1032 => x"4f4d4520",
  1033 => x"53545249",
  1034 => x"4e470000",
  1035 => x"44485259",
  1036 => x"53544f4e",
  1037 => x"45205052",
  1038 => x"4f475241",
  1039 => x"4d2c2031",
  1040 => x"27535420",
  1041 => x"53545249",
  1042 => x"4e470000",
  1043 => x"44687279",
  1044 => x"73746f6e",
  1045 => x"65204265",
  1046 => x"6e63686d",
  1047 => x"61726b2c",
  1048 => x"20566572",
  1049 => x"73696f6e",
  1050 => x"20322e31",
  1051 => x"20284c61",
  1052 => x"6e677561",
  1053 => x"67653a20",
  1054 => x"43290a00",
  1055 => x"50726f67",
  1056 => x"72616d20",
  1057 => x"636f6d70",
  1058 => x"696c6564",
  1059 => x"20776974",
  1060 => x"68202772",
  1061 => x"65676973",
  1062 => x"74657227",
  1063 => x"20617474",
  1064 => x"72696275",
  1065 => x"74650a00",
  1066 => x"45786563",
  1067 => x"7574696f",
  1068 => x"6e207374",
  1069 => x"61727473",
  1070 => x"2c202564",
  1071 => x"2072756e",
  1072 => x"73207468",
  1073 => x"726f7567",
  1074 => x"68204468",
  1075 => x"72797374",
  1076 => x"6f6e650a",
  1077 => x"00000000",
  1078 => x"44485259",
  1079 => x"53544f4e",
  1080 => x"45205052",
  1081 => x"4f475241",
  1082 => x"4d2c2032",
  1083 => x"274e4420",
  1084 => x"53545249",
  1085 => x"4e470000",
  1086 => x"55736572",
  1087 => x"2074696d",
  1088 => x"653a2025",
  1089 => x"640a0000",
  1090 => x"4d696372",
  1091 => x"6f736563",
  1092 => x"6f6e6473",
  1093 => x"20666f72",
  1094 => x"206f6e65",
  1095 => x"2072756e",
  1096 => x"20746872",
  1097 => x"6f756768",
  1098 => x"20446872",
  1099 => x"7973746f",
  1100 => x"6e653a20",
  1101 => x"00000000",
  1102 => x"2564200a",
  1103 => x"00000000",
  1104 => x"44687279",
  1105 => x"73746f6e",
  1106 => x"65732070",
  1107 => x"65722053",
  1108 => x"65636f6e",
  1109 => x"643a2020",
  1110 => x"20202020",
  1111 => x"20202020",
  1112 => x"20202020",
  1113 => x"20202020",
  1114 => x"20202020",
  1115 => x"00000000",
  1116 => x"56415820",
  1117 => x"4d495053",
  1118 => x"20726174",
  1119 => x"696e6720",
  1120 => x"2a203130",
  1121 => x"3030203d",
  1122 => x"20256420",
  1123 => x"0a000000",
  1124 => x"50726f67",
  1125 => x"72616d20",
  1126 => x"636f6d70",
  1127 => x"696c6564",
  1128 => x"20776974",
  1129 => x"686f7574",
  1130 => x"20277265",
  1131 => x"67697374",
  1132 => x"65722720",
  1133 => x"61747472",
  1134 => x"69627574",
  1135 => x"650a0000",
  1136 => x"4d656173",
  1137 => x"75726564",
  1138 => x"2074696d",
  1139 => x"6520746f",
  1140 => x"6f20736d",
  1141 => x"616c6c20",
  1142 => x"746f206f",
  1143 => x"62746169",
  1144 => x"6e206d65",
  1145 => x"616e696e",
  1146 => x"6766756c",
  1147 => x"20726573",
  1148 => x"756c7473",
  1149 => x"0a000000",
  1150 => x"506c6561",
  1151 => x"73652069",
  1152 => x"6e637265",
  1153 => x"61736520",
  1154 => x"6e756d62",
  1155 => x"6572206f",
  1156 => x"66207275",
  1157 => x"6e730a00",
  1158 => x"44485259",
  1159 => x"53544f4e",
  1160 => x"45205052",
  1161 => x"4f475241",
  1162 => x"4d2c2033",
  1163 => x"27524420",
  1164 => x"53545249",
  1165 => x"4e470000",
  1166 => x"000061a8",
  1167 => x"00000000",
	others => x"00000000"
);

begin

process (clk)
begin
	if (clk'event and clk = '1') then
		if (from_zpu.memAWriteEnable = '1') and (from_zpu.memBWriteEnable = '1') and (from_zpu.memAAddr=from_zpu.memBAddr) and (from_zpu.memAWrite/=from_zpu.memBWrite) then
			report "write collision" severity failure;
		end if;
	
		if (from_zpu.memAWriteEnable = '1') then
			ram(to_integer(unsigned(from_zpu.memAAddr(maxAddrBit downto 2)))) := from_zpu.memAWrite;
			to_zpu.memARead <= from_zpu.memAWrite;
		else
			to_zpu.memARead <= ram(to_integer(unsigned(from_zpu.memAAddr(maxAddrBit downto 2))));
		end if;
	end if;
end process;

process (clk)
begin
	if (clk'event and clk = '1') then
		if (from_zpu.memBWriteEnable = '1') then
			ram(to_integer(unsigned(from_zpu.memBAddr(maxAddrBit downto 2)))) := from_zpu.memBWrite;
			to_zpu.memBRead <= from_zpu.memBWrite;
		else
			to_zpu.memBRead <= ram(to_integer(unsigned(from_zpu.memBAddr(maxAddrBit downto 2))));
		end if;
	end if;
end process;


end arch;

