-- ZPU
--
-- Copyright 2004-2008 oharboe - �yvind Harboe - oyvind.harboe@zylin.com
-- Modified by Alastair M. Robinson for the ZPUFlex project.
--
-- The FreeBSD license
-- 
-- Redistribution and use in source and binary forms, with or without
-- modification, are permitted provided that the following conditions
-- are met:
-- 
-- 1. Redistributions of source code must retain the above copyright
--    notice, this list of conditions and the following disclaimer.
-- 2. Redistributions in binary form must reproduce the above
--    copyright notice, this list of conditions and the following
--    disclaimer in the documentation and/or other materials
--    provided with the distribution.
-- 
-- THIS SOFTWARE IS PROVIDED BY THE ZPU PROJECT ``AS IS'' AND ANY
-- EXPRESS OR IMPLIED WARRANTIES, INCLUDING, BUT NOT LIMITED TO,
-- THE IMPLIED WARRANTIES OF MERCHANTABILITY AND FITNESS FOR A
-- PARTICULAR PURPOSE ARE DISCLAIMED. IN NO EVENT SHALL THE
-- ZPU PROJECT OR CONTRIBUTORS BE LIABLE FOR ANY DIRECT,
-- INDIRECT, INCIDENTAL, SPECIAL, EXEMPLARY, OR CONSEQUENTIAL DAMAGES
-- (INCLUDING, BUT NOT LIMITED TO, PROCUREMENT OF SUBSTITUTE GOODS
-- OR SERVICES; LOSS OF USE, DATA, OR PROFITS; OR BUSINESS INTERRUPTION)
-- HOWEVER CAUSED AND ON ANY THEORY OF LIABILITY, WHETHER IN CONTRACT,
-- STRICT LIABILITY, OR TORT (INCLUDING NEGLIGENCE OR OTHERWISE)
-- ARISING IN ANY WAY OUT OF THE USE OF THIS SOFTWARE, EVEN IF
-- ADVISED OF THE POSSIBILITY OF SUCH DAMAGE.
-- 
-- The views and conclusions contained in the software and documentation
-- are those of the authors and should not be interpreted as representing
-- official policies, either expressed or implied, of the ZPU Project.

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;


library work;
use work.zpupkg.all;

entity SDRAMTest_ROM is
generic
	(
		maxAddrBitBRAM : integer := maxAddrBitBRAMLimit -- Specify your actual ROM size to save LEs and unnecessary block RAM usage.
	);
port (
	clk : in std_logic;
	areset : in std_logic := '0';
	from_zpu : in ZPU_ToROM;
	to_zpu : out ZPU_FromROM
);
end SDRAMTest_ROM;

architecture arch of SDRAMTest_ROM is

type ram_type is array(natural range 0 to ((2**(maxAddrBitBRAM+1))/4)-1) of std_logic_vector(wordSize-1 downto 0);

shared variable ram : ram_type :=
(
     0 => x"84808080",
     1 => x"8c0b8480",
     2 => x"8081e004",
     3 => x"00848080",
     4 => x"808c04ff",
     5 => x"0d800404",
     6 => x"40000017",
     7 => x"00000000",
     8 => x"848080a2",
     9 => x"98088480",
    10 => x"80a29c08",
    11 => x"848080a2",
    12 => x"a0088480",
    13 => x"80809808",
    14 => x"2d848080",
    15 => x"a2a00c84",
    16 => x"8080a29c",
    17 => x"0c848080",
    18 => x"a2980c04",
    19 => x"00000000",
    20 => x"00000000",
    21 => x"00000000",
    22 => x"00000000",
    23 => x"00000000",
    24 => x"71fd0608",
    25 => x"72830609",
    26 => x"81058205",
    27 => x"832b2a83",
    28 => x"ffff0652",
    29 => x"0471fc06",
    30 => x"08728306",
    31 => x"09810583",
    32 => x"05101010",
    33 => x"2a81ff06",
    34 => x"520471fd",
    35 => x"060883ff",
    36 => x"ff738306",
    37 => x"09810582",
    38 => x"05832b2b",
    39 => x"09067383",
    40 => x"ffff0673",
    41 => x"83060981",
    42 => x"05820583",
    43 => x"2b0b2b07",
    44 => x"72fc060c",
    45 => x"51510471",
    46 => x"fc060884",
    47 => x"808097cc",
    48 => x"73830610",
    49 => x"10050806",
    50 => x"7381ff06",
    51 => x"73830609",
    52 => x"81058305",
    53 => x"1010102b",
    54 => x"0772fc06",
    55 => x"0c515104",
    56 => x"848080a2",
    57 => x"98708480",
    58 => x"80a3b827",
    59 => x"8e388071",
    60 => x"70840553",
    61 => x"0c848080",
    62 => x"81e50484",
    63 => x"8080808c",
    64 => x"51848080",
    65 => x"92d00402",
    66 => x"c0050d02",
    67 => x"80c4055b",
    68 => x"80707c70",
    69 => x"84055e08",
    70 => x"725f5f5f",
    71 => x"5a7c7084",
    72 => x"055e0857",
    73 => x"80597698",
    74 => x"2a77882b",
    75 => x"58557480",
    76 => x"2e82f338",
    77 => x"7b802e80",
    78 => x"d338805c",
    79 => x"7480e42e",
    80 => x"81de3874",
    81 => x"80f82e81",
    82 => x"d7387480",
    83 => x"e42e81e2",
    84 => x"387480e4",
    85 => x"2680f138",
    86 => x"7480e32e",
    87 => x"80c838a5",
    88 => x"51848080",
    89 => x"868b2d74",
    90 => x"51848080",
    91 => x"868b2d82",
    92 => x"1a811a5a",
    93 => x"5a837925",
    94 => x"ffac3874",
    95 => x"ff9f387e",
    96 => x"848080a2",
    97 => x"980c0280",
    98 => x"c0050d04",
    99 => x"74a52e09",
   100 => x"81069b38",
   101 => x"810b811a",
   102 => x"5a5c8379",
   103 => x"25ff8738",
   104 => x"84808082",
   105 => x"fb047a84",
   106 => x"1c710857",
   107 => x"5c547451",
   108 => x"84808086",
   109 => x"8b2d811a",
   110 => x"811a5a5a",
   111 => x"837925fe",
   112 => x"e5388480",
   113 => x"8082fb04",
   114 => x"7480f32e",
   115 => x"81e53874",
   116 => x"80f82e09",
   117 => x"8106ff87",
   118 => x"387d5380",
   119 => x"58777e24",
   120 => x"82963872",
   121 => x"802e81f9",
   122 => x"38875672",
   123 => x"9c2a7384",
   124 => x"2b545271",
   125 => x"802e8338",
   126 => x"8158b712",
   127 => x"54718924",
   128 => x"8438b012",
   129 => x"547780f0",
   130 => x"38ff1656",
   131 => x"758025db",
   132 => x"38811959",
   133 => x"837925fe",
   134 => x"8d388480",
   135 => x"8082fb04",
   136 => x"7a841c71",
   137 => x"08405c52",
   138 => x"7480e42e",
   139 => x"098106fe",
   140 => x"a0387d54",
   141 => x"8058777e",
   142 => x"24819538",
   143 => x"73802e81",
   144 => x"a0388756",
   145 => x"739c2a74",
   146 => x"842b5552",
   147 => x"71802e83",
   148 => x"388158b7",
   149 => x"12537189",
   150 => x"248438b0",
   151 => x"125377af",
   152 => x"38ff1656",
   153 => x"758025dc",
   154 => x"38811959",
   155 => x"837925fd",
   156 => x"b5388480",
   157 => x"8082fb04",
   158 => x"73518480",
   159 => x"80868b2d",
   160 => x"ff165675",
   161 => x"8025fee3",
   162 => x"38848080",
   163 => x"84910472",
   164 => x"51848080",
   165 => x"868b2dff",
   166 => x"16567580",
   167 => x"25ffa538",
   168 => x"84808084",
   169 => x"e9047984",
   170 => x"8080a298",
   171 => x"0c0280c0",
   172 => x"050d047a",
   173 => x"841c7108",
   174 => x"535c5384",
   175 => x"808086b0",
   176 => x"2d811959",
   177 => x"837925fc",
   178 => x"dd388480",
   179 => x"8082fb04",
   180 => x"ad518480",
   181 => x"80868b2d",
   182 => x"7d098105",
   183 => x"5473fee2",
   184 => x"38b05184",
   185 => x"8080868b",
   186 => x"2d811959",
   187 => x"837925fc",
   188 => x"b5388480",
   189 => x"8082fb04",
   190 => x"ad518480",
   191 => x"80868b2d",
   192 => x"7d098105",
   193 => x"53848080",
   194 => x"83e30402",
   195 => x"f8050d73",
   196 => x"52c00870",
   197 => x"882a7081",
   198 => x"06515151",
   199 => x"70802ef1",
   200 => x"3871c00c",
   201 => x"71848080",
   202 => x"a2980c02",
   203 => x"88050d04",
   204 => x"02e8050d",
   205 => x"80785755",
   206 => x"75708405",
   207 => x"57085380",
   208 => x"5472982a",
   209 => x"73882b54",
   210 => x"5271802e",
   211 => x"a238c008",
   212 => x"70882a70",
   213 => x"81065151",
   214 => x"5170802e",
   215 => x"f13871c0",
   216 => x"0c811581",
   217 => x"15555583",
   218 => x"7425d638",
   219 => x"71ca3874",
   220 => x"848080a2",
   221 => x"980c0298",
   222 => x"050d0402",
   223 => x"f4050d74",
   224 => x"76525380",
   225 => x"71259038",
   226 => x"70527270",
   227 => x"84055408",
   228 => x"ff135351",
   229 => x"71f43802",
   230 => x"8c050d04",
   231 => x"02d4050d",
   232 => x"7c7e5c58",
   233 => x"810b8480",
   234 => x"8097dc58",
   235 => x"5a835976",
   236 => x"08780c77",
   237 => x"08770856",
   238 => x"5473752e",
   239 => x"94387708",
   240 => x"53745284",
   241 => x"808097ec",
   242 => x"51848080",
   243 => x"82872d80",
   244 => x"5a775680",
   245 => x"7b259038",
   246 => x"7a557570",
   247 => x"84055708",
   248 => x"ff165654",
   249 => x"74f43877",
   250 => x"08770856",
   251 => x"5675752e",
   252 => x"94387708",
   253 => x"53745284",
   254 => x"808098ac",
   255 => x"51848080",
   256 => x"82872d80",
   257 => x"5aff1984",
   258 => x"18585978",
   259 => x"8025ff9f",
   260 => x"38798480",
   261 => x"80a2980c",
   262 => x"02ac050d",
   263 => x"0402e405",
   264 => x"0d787a55",
   265 => x"56815785",
   266 => x"aad5aad5",
   267 => x"760cfad5",
   268 => x"aad5aa0b",
   269 => x"8c170ccc",
   270 => x"7634b30b",
   271 => x"8f173475",
   272 => x"085372fc",
   273 => x"e2d5aad5",
   274 => x"2e923875",
   275 => x"08528480",
   276 => x"8098ec51",
   277 => x"84808082",
   278 => x"872d8057",
   279 => x"8c160855",
   280 => x"74fad5aa",
   281 => x"d4b32e93",
   282 => x"388c1608",
   283 => x"52848080",
   284 => x"99a85184",
   285 => x"80808287",
   286 => x"2d805775",
   287 => x"55807425",
   288 => x"8e387470",
   289 => x"84055608",
   290 => x"ff155553",
   291 => x"73f43875",
   292 => x"085473fc",
   293 => x"e2d5aad5",
   294 => x"2e923875",
   295 => x"08528480",
   296 => x"8099e451",
   297 => x"84808082",
   298 => x"872d8057",
   299 => x"8c160853",
   300 => x"72fad5aa",
   301 => x"d4b32e93",
   302 => x"388c1608",
   303 => x"52848080",
   304 => x"9aa05184",
   305 => x"80808287",
   306 => x"2d805776",
   307 => x"848080a2",
   308 => x"980c029c",
   309 => x"050d0402",
   310 => x"e8050d77",
   311 => x"79555680",
   312 => x"c4c4b376",
   313 => x"0c84a2d5",
   314 => x"ccf70b84",
   315 => x"170cf8c4",
   316 => x"e6d5bb0b",
   317 => x"88170cfc",
   318 => x"e6f7ddff",
   319 => x"0b8c170c",
   320 => x"85aad6d5",
   321 => x"aa0b9017",
   322 => x"0c821608",
   323 => x"53728291",
   324 => x"cd88d52e",
   325 => x"8f387252",
   326 => x"8480809a",
   327 => x"dc518480",
   328 => x"8082872d",
   329 => x"86160853",
   330 => x"7286b3de",
   331 => x"91992e8f",
   332 => x"38725284",
   333 => x"80809b98",
   334 => x"51848080",
   335 => x"82872d8a",
   336 => x"16085372",
   337 => x"fad5ef99",
   338 => x"dd2e8f38",
   339 => x"72528480",
   340 => x"809bd451",
   341 => x"84808082",
   342 => x"872d8e16",
   343 => x"085372fe",
   344 => x"f7fdaad5",
   345 => x"2e8f3872",
   346 => x"52848080",
   347 => x"9c905184",
   348 => x"80808287",
   349 => x"2d755580",
   350 => x"74258e38",
   351 => x"74708405",
   352 => x"5608ff15",
   353 => x"555373f4",
   354 => x"38821608",
   355 => x"53728291",
   356 => x"cd88d52e",
   357 => x"8f387252",
   358 => x"8480809c",
   359 => x"cc518480",
   360 => x"8082872d",
   361 => x"86160853",
   362 => x"7286b3de",
   363 => x"91992e8f",
   364 => x"38725284",
   365 => x"80809d88",
   366 => x"51848080",
   367 => x"82872d8a",
   368 => x"16085372",
   369 => x"fad5ef99",
   370 => x"dd2e8f38",
   371 => x"72528480",
   372 => x"809dc451",
   373 => x"84808082",
   374 => x"872d8e16",
   375 => x"085372fe",
   376 => x"f7fdaad5",
   377 => x"2e8f3872",
   378 => x"52848080",
   379 => x"9e805184",
   380 => x"80808287",
   381 => x"2d728480",
   382 => x"80a2980c",
   383 => x"0298050d",
   384 => x"0402cc05",
   385 => x"0d7e5a80",
   386 => x"0b848080",
   387 => x"9ebc5259",
   388 => x"84808082",
   389 => x"872d80e1",
   390 => x"b35780fe",
   391 => x"5dae5184",
   392 => x"8080868b",
   393 => x"2d765c8f",
   394 => x"ffff5876",
   395 => x"bfffff06",
   396 => x"7010101b",
   397 => x"56750c76",
   398 => x"1070962a",
   399 => x"81065657",
   400 => x"74802e85",
   401 => x"38768107",
   402 => x"5776952a",
   403 => x"81065574",
   404 => x"802e8538",
   405 => x"76813257",
   406 => x"ff185877",
   407 => x"8025cc38",
   408 => x"7b578fff",
   409 => x"ff5876bf",
   410 => x"ffff0670",
   411 => x"10101b70",
   412 => x"08575d56",
   413 => x"74762e81",
   414 => x"8b388079",
   415 => x"53848080",
   416 => x"9ecc525b",
   417 => x"84808082",
   418 => x"872d7454",
   419 => x"75537552",
   420 => x"8480809e",
   421 => x"e0518480",
   422 => x"8082872d",
   423 => x"7a597610",
   424 => x"70962a81",
   425 => x"06565774",
   426 => x"802e8538",
   427 => x"76810757",
   428 => x"76952a81",
   429 => x"065c7b80",
   430 => x"2e853876",
   431 => x"813257ff",
   432 => x"18587780",
   433 => x"25ff9f38",
   434 => x"76107096",
   435 => x"2a810659",
   436 => x"5777802e",
   437 => x"85387681",
   438 => x"07577695",
   439 => x"2a81065c",
   440 => x"7b802e85",
   441 => x"38768132",
   442 => x"57ff1d5d",
   443 => x"7cfeae38",
   444 => x"8a518480",
   445 => x"80868b2d",
   446 => x"7a848080",
   447 => x"a2980c02",
   448 => x"b4050d04",
   449 => x"81195984",
   450 => x"80808d9e",
   451 => x"0402c805",
   452 => x"0d7f5d80",
   453 => x"61922bff",
   454 => x"055b5b80",
   455 => x"e1b30b84",
   456 => x"80809f88",
   457 => x"52578480",
   458 => x"8082872d",
   459 => x"7a7a2781",
   460 => x"9e387c7a",
   461 => x"5a587678",
   462 => x"0c761070",
   463 => x"962a7081",
   464 => x"06515757",
   465 => x"75802e85",
   466 => x"38768107",
   467 => x"5776952a",
   468 => x"70810651",
   469 => x"5675802e",
   470 => x"85387681",
   471 => x"3257ff19",
   472 => x"84195959",
   473 => x"78d03880",
   474 => x"e1b35780",
   475 => x"7a2780df",
   476 => x"387c5877",
   477 => x"08567577",
   478 => x"2e80e838",
   479 => x"807b5384",
   480 => x"80809ecc",
   481 => x"525c8480",
   482 => x"8082872d",
   483 => x"7d557554",
   484 => x"76537852",
   485 => x"8480809f",
   486 => x"9c518480",
   487 => x"8082872d",
   488 => x"7b5b7610",
   489 => x"70962a81",
   490 => x"065e577c",
   491 => x"802e8538",
   492 => x"76810757",
   493 => x"76952a81",
   494 => x"065d7c80",
   495 => x"2e853876",
   496 => x"81325781",
   497 => x"19841959",
   498 => x"59797926",
   499 => x"ffa5388a",
   500 => x"51848080",
   501 => x"868b2d7b",
   502 => x"848080a2",
   503 => x"980c02b8",
   504 => x"050d0481",
   505 => x"1b5b8480",
   506 => x"808fa204",
   507 => x"02cc050d",
   508 => x"7e605e58",
   509 => x"815a805b",
   510 => x"80c07a58",
   511 => x"5c85ada9",
   512 => x"89bb780c",
   513 => x"79598156",
   514 => x"97557676",
   515 => x"07822b78",
   516 => x"11515485",
   517 => x"ada989bb",
   518 => x"740c7510",
   519 => x"ff165656",
   520 => x"748025e6",
   521 => x"38761081",
   522 => x"1a5a5798",
   523 => x"7925d738",
   524 => x"7756807d",
   525 => x"2590387c",
   526 => x"55757084",
   527 => x"055708ff",
   528 => x"16565474",
   529 => x"f4388157",
   530 => x"ff8787a5",
   531 => x"c3780c97",
   532 => x"5976822b",
   533 => x"78117008",
   534 => x"5f56567c",
   535 => x"ff8787a5",
   536 => x"c32e80cc",
   537 => x"38740854",
   538 => x"7385ada9",
   539 => x"89bb2e94",
   540 => x"38807508",
   541 => x"54765384",
   542 => x"80809fd0",
   543 => x"525a8480",
   544 => x"8082872d",
   545 => x"7610ff1a",
   546 => x"5a577880",
   547 => x"25c3387a",
   548 => x"822b5675",
   549 => x"b1387b52",
   550 => x"8480809f",
   551 => x"f0518480",
   552 => x"8082872d",
   553 => x"7b848080",
   554 => x"a2980c02",
   555 => x"b4050d04",
   556 => x"7a770777",
   557 => x"10ff1b5b",
   558 => x"585b7880",
   559 => x"25ff9238",
   560 => x"84808091",
   561 => x"8f047552",
   562 => x"848080a0",
   563 => x"ac518480",
   564 => x"8082872d",
   565 => x"75992a81",
   566 => x"32810670",
   567 => x"09810571",
   568 => x"07700970",
   569 => x"9f2c7d06",
   570 => x"79109fff",
   571 => x"fffc0660",
   572 => x"812a415a",
   573 => x"5d575859",
   574 => x"75da3879",
   575 => x"09810570",
   576 => x"7b079f2a",
   577 => x"55567bbf",
   578 => x"26843873",
   579 => x"9d388170",
   580 => x"53848080",
   581 => x"9ff0525c",
   582 => x"84808082",
   583 => x"872d7b84",
   584 => x"8080a298",
   585 => x"0c02b405",
   586 => x"0d048480",
   587 => x"80a0c451",
   588 => x"84808082",
   589 => x"872d7b52",
   590 => x"8480809f",
   591 => x"f0518480",
   592 => x"8082872d",
   593 => x"7b848080",
   594 => x"a2980c02",
   595 => x"b4050d04",
   596 => x"02cc050d",
   597 => x"810b8480",
   598 => x"8097dc5a",
   599 => x"5a835b78",
   600 => x"08800c80",
   601 => x"08790858",
   602 => x"5675772e",
   603 => x"94388008",
   604 => x"53765284",
   605 => x"808097ec",
   606 => x"51848080",
   607 => x"82872d80",
   608 => x"5a807059",
   609 => x"57777084",
   610 => x"05590881",
   611 => x"185856a0",
   612 => x"807724f1",
   613 => x"38800879",
   614 => x"08585877",
   615 => x"772e9438",
   616 => x"80085376",
   617 => x"52848080",
   618 => x"98ac5184",
   619 => x"80808287",
   620 => x"2d805aff",
   621 => x"1b841a5a",
   622 => x"5b7a8025",
   623 => x"ffa13879",
   624 => x"802e8d38",
   625 => x"848080a1",
   626 => x"90518480",
   627 => x"8082872d",
   628 => x"815985aa",
   629 => x"d5aad50b",
   630 => x"800cfad5",
   631 => x"aad5aa0b",
   632 => x"8c0ccc0b",
   633 => x"8034b30b",
   634 => x"8f348008",
   635 => x"5776fce2",
   636 => x"d5aad52e",
   637 => x"92388008",
   638 => x"52848080",
   639 => x"98ec5184",
   640 => x"80808287",
   641 => x"2d80598c",
   642 => x"085a79fa",
   643 => x"d5aad4b3",
   644 => x"2e92388c",
   645 => x"08528480",
   646 => x"8099a851",
   647 => x"84808082",
   648 => x"872d8059",
   649 => x"80705957",
   650 => x"77708405",
   651 => x"59088118",
   652 => x"5856a080",
   653 => x"7724f138",
   654 => x"80085b7a",
   655 => x"fce2d5aa",
   656 => x"d52e9238",
   657 => x"80085284",
   658 => x"808099e4",
   659 => x"51848080",
   660 => x"82872d80",
   661 => x"598c0856",
   662 => x"75fad5aa",
   663 => x"d4b32e82",
   664 => x"d0388c08",
   665 => x"52848080",
   666 => x"9aa05184",
   667 => x"80808287",
   668 => x"2da08052",
   669 => x"80518480",
   670 => x"808fec2d",
   671 => x"848080a2",
   672 => x"98085a84",
   673 => x"8080a298",
   674 => x"08802e8d",
   675 => x"38848080",
   676 => x"a1b45184",
   677 => x"80808287",
   678 => x"2d807a90",
   679 => x"808029ff",
   680 => x"055a5b80",
   681 => x"e1b30b84",
   682 => x"80809f88",
   683 => x"52578480",
   684 => x"8082872d",
   685 => x"7a587a79",
   686 => x"2781a238",
   687 => x"77822b77",
   688 => x"710c5676",
   689 => x"1070962a",
   690 => x"70810651",
   691 => x"57577580",
   692 => x"2e853876",
   693 => x"81075776",
   694 => x"952a7081",
   695 => x"06515675",
   696 => x"802e8538",
   697 => x"76813257",
   698 => x"81185878",
   699 => x"7826cd38",
   700 => x"80e1b357",
   701 => x"80587779",
   702 => x"2780e238",
   703 => x"77822b70",
   704 => x"08515675",
   705 => x"772e81a0",
   706 => x"38807b53",
   707 => x"8480809e",
   708 => x"cc525c84",
   709 => x"80808287",
   710 => x"2d7c5575",
   711 => x"54765377",
   712 => x"52848080",
   713 => x"9f9c5184",
   714 => x"80808287",
   715 => x"2d7b5b76",
   716 => x"1070962a",
   717 => x"70810651",
   718 => x"57577580",
   719 => x"2e853876",
   720 => x"81075776",
   721 => x"952a7081",
   722 => x"06515675",
   723 => x"802e8538",
   724 => x"76813257",
   725 => x"81185878",
   726 => x"7826ffa0",
   727 => x"388a5184",
   728 => x"8080868b",
   729 => x"2d7b802e",
   730 => x"8d388480",
   731 => x"80a1cc51",
   732 => x"84808082",
   733 => x"872d7952",
   734 => x"80518480",
   735 => x"808c812d",
   736 => x"848080a2",
   737 => x"9808802e",
   738 => x"fbca3884",
   739 => x"8080a1e4",
   740 => x"51848080",
   741 => x"82872d81",
   742 => x"0b848080",
   743 => x"97dc5a5a",
   744 => x"835b8480",
   745 => x"8092df04",
   746 => x"811b5b84",
   747 => x"808096af",
   748 => x"0478802e",
   749 => x"fdbb3884",
   750 => x"8080a1fc",
   751 => x"51848080",
   752 => x"82872d84",
   753 => x"808094f1",
   754 => x"04000000",
   755 => x"00ffffff",
   756 => x"ff00ffff",
   757 => x"ffff00ff",
   758 => x"ffffff00",
   759 => x"00000000",
   760 => x"55555555",
   761 => x"aaaaaaaa",
   762 => x"ffffffff",
   763 => x"53616e69",
   764 => x"74792063",
   765 => x"6865636b",
   766 => x"20666169",
   767 => x"6c656420",
   768 => x"28626566",
   769 => x"6f726520",
   770 => x"63616368",
   771 => x"65207265",
   772 => x"66726573",
   773 => x"6829206f",
   774 => x"6e203078",
   775 => x"25642028",
   776 => x"676f7420",
   777 => x"30782564",
   778 => x"290a0000",
   779 => x"53616e69",
   780 => x"74792063",
   781 => x"6865636b",
   782 => x"20666169",
   783 => x"6c656420",
   784 => x"28616674",
   785 => x"65722063",
   786 => x"61636865",
   787 => x"20726566",
   788 => x"72657368",
   789 => x"29206f6e",
   790 => x"20307825",
   791 => x"64202867",
   792 => x"6f742030",
   793 => x"78256429",
   794 => x"0a000000",
   795 => x"42797465",
   796 => x"20636865",
   797 => x"636b2066",
   798 => x"61696c65",
   799 => x"64202862",
   800 => x"65666f72",
   801 => x"65206361",
   802 => x"63686520",
   803 => x"72656672",
   804 => x"65736829",
   805 => x"20617420",
   806 => x"30202867",
   807 => x"6f742030",
   808 => x"78256429",
   809 => x"0a000000",
   810 => x"42797465",
   811 => x"20636865",
   812 => x"636b2066",
   813 => x"61696c65",
   814 => x"64202862",
   815 => x"65666f72",
   816 => x"65206361",
   817 => x"63686520",
   818 => x"72656672",
   819 => x"65736829",
   820 => x"20617420",
   821 => x"33202867",
   822 => x"6f742030",
   823 => x"78256429",
   824 => x"0a000000",
   825 => x"42797465",
   826 => x"20636865",
   827 => x"636b2066",
   828 => x"61696c65",
   829 => x"64202861",
   830 => x"66746572",
   831 => x"20636163",
   832 => x"68652072",
   833 => x"65667265",
   834 => x"73682920",
   835 => x"61742030",
   836 => x"2028676f",
   837 => x"74203078",
   838 => x"2564290a",
   839 => x"00000000",
   840 => x"42797465",
   841 => x"20636865",
   842 => x"636b2066",
   843 => x"61696c65",
   844 => x"64202861",
   845 => x"66746572",
   846 => x"20636163",
   847 => x"68652072",
   848 => x"65667265",
   849 => x"73682920",
   850 => x"61742033",
   851 => x"2028676f",
   852 => x"74203078",
   853 => x"2564290a",
   854 => x"00000000",
   855 => x"416c6967",
   856 => x"6e206368",
   857 => x"65636b20",
   858 => x"6661696c",
   859 => x"65642028",
   860 => x"6265666f",
   861 => x"72652063",
   862 => x"61636865",
   863 => x"20726566",
   864 => x"72657368",
   865 => x"29206174",
   866 => x"20322028",
   867 => x"676f7420",
   868 => x"30782564",
   869 => x"290a0000",
   870 => x"416c6967",
   871 => x"6e206368",
   872 => x"65636b20",
   873 => x"6661696c",
   874 => x"65642028",
   875 => x"6265666f",
   876 => x"72652063",
   877 => x"61636865",
   878 => x"20726566",
   879 => x"72657368",
   880 => x"29206174",
   881 => x"20362028",
   882 => x"676f7420",
   883 => x"30782564",
   884 => x"290a0000",
   885 => x"416c6967",
   886 => x"6e206368",
   887 => x"65636b20",
   888 => x"6661696c",
   889 => x"65642028",
   890 => x"6265666f",
   891 => x"72652063",
   892 => x"61636865",
   893 => x"20726566",
   894 => x"72657368",
   895 => x"29206174",
   896 => x"20313020",
   897 => x"28676f74",
   898 => x"20307825",
   899 => x"64290a00",
   900 => x"416c6967",
   901 => x"6e206368",
   902 => x"65636b20",
   903 => x"6661696c",
   904 => x"65642028",
   905 => x"6265666f",
   906 => x"72652063",
   907 => x"61636865",
   908 => x"20726566",
   909 => x"72657368",
   910 => x"29206174",
   911 => x"20313420",
   912 => x"28676f74",
   913 => x"20307825",
   914 => x"64290a00",
   915 => x"416c6967",
   916 => x"6e206368",
   917 => x"65636b20",
   918 => x"6661696c",
   919 => x"65642028",
   920 => x"61667465",
   921 => x"72206361",
   922 => x"63686520",
   923 => x"72656672",
   924 => x"65736829",
   925 => x"20617420",
   926 => x"32202867",
   927 => x"6f742030",
   928 => x"78256429",
   929 => x"0a000000",
   930 => x"416c6967",
   931 => x"6e206368",
   932 => x"65636b20",
   933 => x"6661696c",
   934 => x"65642028",
   935 => x"61667465",
   936 => x"72206361",
   937 => x"63686520",
   938 => x"72656672",
   939 => x"65736829",
   940 => x"20617420",
   941 => x"36202867",
   942 => x"6f742030",
   943 => x"78256429",
   944 => x"0a000000",
   945 => x"416c6967",
   946 => x"6e206368",
   947 => x"65636b20",
   948 => x"6661696c",
   949 => x"65642028",
   950 => x"61667465",
   951 => x"72206361",
   952 => x"63686520",
   953 => x"72656672",
   954 => x"65736829",
   955 => x"20617420",
   956 => x"31302028",
   957 => x"676f7420",
   958 => x"30782564",
   959 => x"290a0000",
   960 => x"416c6967",
   961 => x"6e206368",
   962 => x"65636b20",
   963 => x"6661696c",
   964 => x"65642028",
   965 => x"61667465",
   966 => x"72206361",
   967 => x"63686520",
   968 => x"72656672",
   969 => x"65736829",
   970 => x"20617420",
   971 => x"31342028",
   972 => x"676f7420",
   973 => x"30782564",
   974 => x"290a0000",
   975 => x"43686563",
   976 => x"6b696e67",
   977 => x"206d656d",
   978 => x"6f727900",
   979 => x"30782564",
   980 => x"20676f6f",
   981 => x"64207265",
   982 => x"6164732c",
   983 => x"20000000",
   984 => x"4572726f",
   985 => x"72206174",
   986 => x"20307825",
   987 => x"642c2065",
   988 => x"78706563",
   989 => x"74656420",
   990 => x"30782564",
   991 => x"2c20676f",
   992 => x"74203078",
   993 => x"25640a00",
   994 => x"4c696e65",
   995 => x"6172206d",
   996 => x"656d6f72",
   997 => x"79206368",
   998 => x"65636b00",
   999 => x"4572726f",
  1000 => x"72206174",
  1001 => x"20307825",
  1002 => x"642c2065",
  1003 => x"78706563",
  1004 => x"74656420",
  1005 => x"30782564",
  1006 => x"2c20676f",
  1007 => x"74203078",
  1008 => x"2564206f",
  1009 => x"6e20726f",
  1010 => x"756e6420",
  1011 => x"25640a00",
  1012 => x"42616420",
  1013 => x"64617461",
  1014 => x"20666f75",
  1015 => x"6e642061",
  1016 => x"74203078",
  1017 => x"25642028",
  1018 => x"30782564",
  1019 => x"290a0000",
  1020 => x"53445241",
  1021 => x"4d207369",
  1022 => x"7a652028",
  1023 => x"61737375",
  1024 => x"6d696e67",
  1025 => x"206e6f20",
  1026 => x"61646472",
  1027 => x"65737320",
  1028 => x"6661756c",
  1029 => x"74732920",
  1030 => x"69732030",
  1031 => x"78256420",
  1032 => x"6d656761",
  1033 => x"62797465",
  1034 => x"730a0000",
  1035 => x"416c6961",
  1036 => x"73657320",
  1037 => x"666f756e",
  1038 => x"64206174",
  1039 => x"20307825",
  1040 => x"640a0000",
  1041 => x"28416c69",
  1042 => x"61736573",
  1043 => x"2070726f",
  1044 => x"6261626c",
  1045 => x"79207369",
  1046 => x"6d706c79",
  1047 => x"20696e64",
  1048 => x"69636174",
  1049 => x"65207468",
  1050 => x"61742052",
  1051 => x"414d0a69",
  1052 => x"7320736d",
  1053 => x"616c6c65",
  1054 => x"72207468",
  1055 => x"616e2036",
  1056 => x"34206d65",
  1057 => x"67616279",
  1058 => x"74657329",
  1059 => x"0a000000",
  1060 => x"46697273",
  1061 => x"74207374",
  1062 => x"61676520",
  1063 => x"73616e69",
  1064 => x"74792063",
  1065 => x"6865636b",
  1066 => x"20706173",
  1067 => x"7365642e",
  1068 => x"0a000000",
  1069 => x"41646472",
  1070 => x"65737320",
  1071 => x"63686563",
  1072 => x"6b207061",
  1073 => x"73736564",
  1074 => x"2e0a0000",
  1075 => x"4c696e65",
  1076 => x"61722063",
  1077 => x"6865636b",
  1078 => x"20706173",
  1079 => x"7365642e",
  1080 => x"0a0a0000",
  1081 => x"4c465352",
  1082 => x"20636865",
  1083 => x"636b2070",
  1084 => x"61737365",
  1085 => x"642e0a0a",
  1086 => x"00000000",
  1087 => x"42797465",
  1088 => x"20286471",
  1089 => x"6d292063",
  1090 => x"6865636b",
  1091 => x"20706173",
  1092 => x"7365640a",
  1093 => x"00000000",
	others => x"00000000"
);

begin

process (clk)
begin
	if (clk'event and clk = '1') then
		if (from_zpu.memAWriteEnable = '1') and (from_zpu.memBWriteEnable = '1') and (from_zpu.memAAddr=from_zpu.memBAddr) and (from_zpu.memAWrite/=from_zpu.memBWrite) then
			report "write collision" severity failure;
		end if;
	
		if (from_zpu.memAWriteEnable = '1') then
			ram(to_integer(unsigned(from_zpu.memAAddr(maxAddrBitBRAM downto 2)))) := from_zpu.memAWrite;
			to_zpu.memARead <= from_zpu.memAWrite;
		else
			to_zpu.memARead <= ram(to_integer(unsigned(from_zpu.memAAddr(maxAddrBitBRAM downto 2))));
		end if;
	end if;
end process;

process (clk)
begin
	if (clk'event and clk = '1') then
		if (from_zpu.memBWriteEnable = '1') then
			ram(to_integer(unsigned(from_zpu.memBAddr(maxAddrBitBRAM downto 2)))) := from_zpu.memBWrite;
			to_zpu.memBRead <= from_zpu.memBWrite;
		else
			to_zpu.memBRead <= ram(to_integer(unsigned(from_zpu.memBAddr(maxAddrBitBRAM downto 2))));
		end if;
	end if;
end process;


end arch;

