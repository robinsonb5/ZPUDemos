-- ZPU
--
-- Copyright 2004-2008 oharboe - �yvind Harboe - oyvind.harboe@zylin.com
-- Modified by Alastair M. Robinson for the ZPUFlex project.
--
-- The FreeBSD license
-- 
-- Redistribution and use in source and binary forms, with or without
-- modification, are permitted provided that the following conditions
-- are met:
-- 
-- 1. Redistributions of source code must retain the above copyright
--    notice, this list of conditions and the following disclaimer.
-- 2. Redistributions in binary form must reproduce the above
--    copyright notice, this list of conditions and the following
--    disclaimer in the documentation and/or other materials
--    provided with the distribution.
-- 
-- THIS SOFTWARE IS PROVIDED BY THE ZPU PROJECT ``AS IS'' AND ANY
-- EXPRESS OR IMPLIED WARRANTIES, INCLUDING, BUT NOT LIMITED TO,
-- THE IMPLIED WARRANTIES OF MERCHANTABILITY AND FITNESS FOR A
-- PARTICULAR PURPOSE ARE DISCLAIMED. IN NO EVENT SHALL THE
-- ZPU PROJECT OR CONTRIBUTORS BE LIABLE FOR ANY DIRECT,
-- INDIRECT, INCIDENTAL, SPECIAL, EXEMPLARY, OR CONSEQUENTIAL DAMAGES
-- (INCLUDING, BUT NOT LIMITED TO, PROCUREMENT OF SUBSTITUTE GOODS
-- OR SERVICES; LOSS OF USE, DATA, OR PROFITS; OR BUSINESS INTERRUPTION)
-- HOWEVER CAUSED AND ON ANY THEORY OF LIABILITY, WHETHER IN CONTRACT,
-- STRICT LIABILITY, OR TORT (INCLUDING NEGLIGENCE OR OTHERWISE)
-- ARISING IN ANY WAY OUT OF THE USE OF THIS SOFTWARE, EVEN IF
-- ADVISED OF THE POSSIBILITY OF SUCH DAMAGE.
-- 
-- The views and conclusions contained in the software and documentation
-- are those of the authors and should not be interpreted as representing
-- official policies, either expressed or implied, of the ZPU Project.

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;


library work;
use work.zpu_config.all;
use work.zpupkg.all;

entity SDRAMTest_ROM is
generic
	(
		maxAddrBit : integer := maxAddrBitBRAMLimit -- Specify your actual ROM size to save LEs and unnecessary block RAM usage.
	);
port (
	clk : in std_logic;
	areset : in std_logic := '0';
	from_zpu : in ZPU_ToROM;
	to_zpu : out ZPU_FromROM
);
end SDRAMTest_ROM;

architecture arch of SDRAMTest_ROM is

type ram_type is array(natural range 0 to ((2**(maxAddrBit+1))/4)-1) of std_logic_vector(wordSize-1 downto 0);

shared variable ram : ram_type :=
(
     0 => x"0ba08080",
     1 => x"e2040000",
     2 => x"8004a080",
     3 => x"808a0471",
     4 => x"fd060872",
     5 => x"83060981",
     6 => x"05820583",
     7 => x"2b2a83ff",
     8 => x"ff065204",
     9 => x"71fc0608",
    10 => x"72830609",
    11 => x"81058305",
    12 => x"1010102a",
    13 => x"81ff0652",
    14 => x"0471fc06",
    15 => x"080ba080",
    16 => x"93847383",
    17 => x"06101005",
    18 => x"08067381",
    19 => x"ff067383",
    20 => x"06098105",
    21 => x"83051010",
    22 => x"102b0772",
    23 => x"fc060c51",
    24 => x"5104a080",
    25 => x"808a0ba0",
    26 => x"808cd704",
    27 => x"0002c005",
    28 => x"0d0280c4",
    29 => x"05a0809a",
    30 => x"845a5c80",
    31 => x"7c708405",
    32 => x"5e08715f",
    33 => x"5f577d70",
    34 => x"84055f08",
    35 => x"56805875",
    36 => x"982a7688",
    37 => x"2b575574",
    38 => x"802e8384",
    39 => x"387c802e",
    40 => x"80c23880",
    41 => x"5d7480e4",
    42 => x"2e81b638",
    43 => x"7480e426",
    44 => x"80eb3874",
    45 => x"80e32e80",
    46 => x"c438a551",
    47 => x"a08084ac",
    48 => x"2d7451a0",
    49 => x"8084ac2d",
    50 => x"82175781",
    51 => x"18588378",
    52 => x"25ffbc38",
    53 => x"74ffaf38",
    54 => x"7ea08099",
    55 => x"a40c0280",
    56 => x"c0050d04",
    57 => x"74a52e09",
    58 => x"81069a38",
    59 => x"810b8119",
    60 => x"595d8378",
    61 => x"25ff9838",
    62 => x"a08081d4",
    63 => x"047b841d",
    64 => x"7108575d",
    65 => x"5a7451a0",
    66 => x"8084ac2d",
    67 => x"81178119",
    68 => x"59578378",
    69 => x"25fef838",
    70 => x"a08081d4",
    71 => x"047480f3",
    72 => x"2e098106",
    73 => x"ff94387b",
    74 => x"841d7108",
    75 => x"70545b5d",
    76 => x"54a08084",
    77 => x"d22d800b",
    78 => x"ff115553",
    79 => x"807325ff",
    80 => x"8a387870",
    81 => x"81055aa0",
    82 => x"8080a42d",
    83 => x"705255a0",
    84 => x"8084ac2d",
    85 => x"811774ff",
    86 => x"16565457",
    87 => x"a08082bc",
    88 => x"047b841d",
    89 => x"7108a080",
    90 => x"9a840ba0",
    91 => x"8099b461",
    92 => x"5f585e52",
    93 => x"5d537280",
    94 => x"c238b00b",
    95 => x"a08099b4",
    96 => x"0ba08080",
    97 => x"b92d8114",
    98 => x"54ff1454",
    99 => x"73a08080",
   100 => x"a42d7b70",
   101 => x"81055da0",
   102 => x"8080b92d",
   103 => x"811a5a73",
   104 => x"a08099b4",
   105 => x"2e098106",
   106 => x"e038807b",
   107 => x"a08080b9",
   108 => x"2d79ff11",
   109 => x"5553a080",
   110 => x"82bc048a",
   111 => x"527251a0",
   112 => x"8090972d",
   113 => x"a08099a4",
   114 => x"08a08093",
   115 => x"9405a080",
   116 => x"80a42d74",
   117 => x"70810556",
   118 => x"a08080b9",
   119 => x"2d8a5272",
   120 => x"51a0808f",
   121 => x"dd2da080",
   122 => x"99a40853",
   123 => x"a08099a4",
   124 => x"08c93873",
   125 => x"a08099b4",
   126 => x"2effaf38",
   127 => x"ff145473",
   128 => x"a08080a4",
   129 => x"2d7b7081",
   130 => x"055da080",
   131 => x"80b92d81",
   132 => x"1a5a73a0",
   133 => x"8099b42e",
   134 => x"ff9038a0",
   135 => x"80838904",
   136 => x"76a08099",
   137 => x"a40c0280",
   138 => x"c0050d04",
   139 => x"02f8050d",
   140 => x"7352ff84",
   141 => x"0870882a",
   142 => x"70810651",
   143 => x"51517080",
   144 => x"2ef03871",
   145 => x"ff840c71",
   146 => x"a08099a4",
   147 => x"0c028805",
   148 => x"0d0402f0",
   149 => x"050d7553",
   150 => x"8073a080",
   151 => x"80a42d52",
   152 => x"5470742e",
   153 => x"a8387052",
   154 => x"811353ff",
   155 => x"84087088",
   156 => x"2a708106",
   157 => x"51515170",
   158 => x"802ef038",
   159 => x"71ff840c",
   160 => x"811473a0",
   161 => x"8080a42d",
   162 => x"535471dc",
   163 => x"3873a080",
   164 => x"99a40c02",
   165 => x"90050d04",
   166 => x"02f4050d",
   167 => x"74765253",
   168 => x"80712590",
   169 => x"38705272",
   170 => x"70840554",
   171 => x"08ff1353",
   172 => x"5171f438",
   173 => x"028c050d",
   174 => x"0402d405",
   175 => x"0d7c7e5c",
   176 => x"58810ba0",
   177 => x"8093a858",
   178 => x"5a835976",
   179 => x"08780c77",
   180 => x"08770856",
   181 => x"5473752e",
   182 => x"92387708",
   183 => x"537452a0",
   184 => x"8093b851",
   185 => x"a08080ed",
   186 => x"2d805a77",
   187 => x"56807b25",
   188 => x"90387a55",
   189 => x"75708405",
   190 => x"5708ff16",
   191 => x"565474f4",
   192 => x"38770877",
   193 => x"08565675",
   194 => x"752e9238",
   195 => x"77085374",
   196 => x"52a08093",
   197 => x"f851a080",
   198 => x"80ed2d80",
   199 => x"5aff1984",
   200 => x"18585978",
   201 => x"8025ffa3",
   202 => x"3879a080",
   203 => x"99a40c02",
   204 => x"ac050d04",
   205 => x"02e4050d",
   206 => x"787a5556",
   207 => x"815785aa",
   208 => x"d5aad576",
   209 => x"0cfad5aa",
   210 => x"d5aa0b8c",
   211 => x"170ccc76",
   212 => x"a08080b9",
   213 => x"2db30b8f",
   214 => x"17a08080",
   215 => x"b92d7508",
   216 => x"5372fce2",
   217 => x"d5aad52e",
   218 => x"90387508",
   219 => x"52a08094",
   220 => x"b851a080",
   221 => x"80ed2d80",
   222 => x"578c1608",
   223 => x"5574fad5",
   224 => x"aad4b32e",
   225 => x"91388c16",
   226 => x"0852a080",
   227 => x"94f451a0",
   228 => x"8080ed2d",
   229 => x"80577555",
   230 => x"8074258e",
   231 => x"38747084",
   232 => x"055608ff",
   233 => x"15555373",
   234 => x"f4387508",
   235 => x"5473fce2",
   236 => x"d5aad52e",
   237 => x"90387508",
   238 => x"52a08095",
   239 => x"b051a080",
   240 => x"80ed2d80",
   241 => x"578c1608",
   242 => x"5372fad5",
   243 => x"aad4b32e",
   244 => x"91388c16",
   245 => x"0852a080",
   246 => x"95ec51a0",
   247 => x"8080ed2d",
   248 => x"805776a0",
   249 => x"8099a40c",
   250 => x"029c050d",
   251 => x"0402c405",
   252 => x"0d605b80",
   253 => x"62908080",
   254 => x"29ff05a0",
   255 => x"8096a853",
   256 => x"405aa080",
   257 => x"80ed2d80",
   258 => x"e1b35780",
   259 => x"fe5eae51",
   260 => x"a08084ac",
   261 => x"2d761070",
   262 => x"962a8106",
   263 => x"56577480",
   264 => x"2e853876",
   265 => x"81075776",
   266 => x"952a8106",
   267 => x"5877802e",
   268 => x"85387681",
   269 => x"32577877",
   270 => x"077f0677",
   271 => x"5e598fff",
   272 => x"ff5876bf",
   273 => x"ffff0670",
   274 => x"7a32822b",
   275 => x"7c115157",
   276 => x"760c7610",
   277 => x"70962a81",
   278 => x"06565774",
   279 => x"802e8538",
   280 => x"76810757",
   281 => x"76952a81",
   282 => x"06557480",
   283 => x"2e853876",
   284 => x"813257ff",
   285 => x"18587780",
   286 => x"25c8387c",
   287 => x"578fffff",
   288 => x"5876bfff",
   289 => x"ff06707a",
   290 => x"32822b7c",
   291 => x"05700857",
   292 => x"5e567476",
   293 => x"2e80e438",
   294 => x"807a53a0",
   295 => x"8096b852",
   296 => x"5ca08080",
   297 => x"ed2d7454",
   298 => x"75537552",
   299 => x"a08096cc",
   300 => x"51a08080",
   301 => x"ed2d7b5a",
   302 => x"76107096",
   303 => x"2a810657",
   304 => x"5775802e",
   305 => x"85387681",
   306 => x"07577695",
   307 => x"2a810655",
   308 => x"74802e85",
   309 => x"38768132",
   310 => x"57ff1858",
   311 => x"778025ff",
   312 => x"a038ff1e",
   313 => x"5e7dfea6",
   314 => x"388a51a0",
   315 => x"8084ac2d",
   316 => x"7ba08099",
   317 => x"a40c02bc",
   318 => x"050d0481",
   319 => x"1a5aa080",
   320 => x"89b80402",
   321 => x"cc050d7e",
   322 => x"605e5881",
   323 => x"5a805b80",
   324 => x"c07a585c",
   325 => x"85ada989",
   326 => x"bb780c79",
   327 => x"59815697",
   328 => x"55767607",
   329 => x"822b7811",
   330 => x"515485ad",
   331 => x"a989bb74",
   332 => x"0c7510ff",
   333 => x"16565674",
   334 => x"8025e638",
   335 => x"7610811a",
   336 => x"5a579879",
   337 => x"25d73877",
   338 => x"56807d25",
   339 => x"90387c55",
   340 => x"75708405",
   341 => x"5708ff16",
   342 => x"565474f4",
   343 => x"388157ff",
   344 => x"8787a5c3",
   345 => x"780c9759",
   346 => x"76822b78",
   347 => x"1170085f",
   348 => x"56567cff",
   349 => x"8787a5c3",
   350 => x"2e80c738",
   351 => x"74085473",
   352 => x"85ada989",
   353 => x"bb2e9238",
   354 => x"80750854",
   355 => x"7653a080",
   356 => x"96f4525a",
   357 => x"a08080ed",
   358 => x"2d7610ff",
   359 => x"1a5a5778",
   360 => x"8025c538",
   361 => x"7a822b56",
   362 => x"75ad387b",
   363 => x"52a08097",
   364 => x"9451a080",
   365 => x"80ed2d7b",
   366 => x"a08099a4",
   367 => x"0c02b405",
   368 => x"0d047a77",
   369 => x"077710ff",
   370 => x"1b5b585b",
   371 => x"788025ff",
   372 => x"9738a080",
   373 => x"8ba40475",
   374 => x"52a08097",
   375 => x"d051a080",
   376 => x"80ed2d75",
   377 => x"992a8132",
   378 => x"81067009",
   379 => x"81057107",
   380 => x"7009709f",
   381 => x"2c7d0679",
   382 => x"109fffff",
   383 => x"fc066081",
   384 => x"2a415a5d",
   385 => x"57585975",
   386 => x"da387909",
   387 => x"8105707b",
   388 => x"079f2a55",
   389 => x"567bbf26",
   390 => x"8438739a",
   391 => x"38817053",
   392 => x"a0809794",
   393 => x"525ca080",
   394 => x"80ed2d7b",
   395 => x"a08099a4",
   396 => x"0c02b405",
   397 => x"0d04a080",
   398 => x"97e851a0",
   399 => x"8080ed2d",
   400 => x"7b52a080",
   401 => x"979451a0",
   402 => x"8080ed2d",
   403 => x"7ba08099",
   404 => x"a40c02b4",
   405 => x"050d0402",
   406 => x"dc050d88",
   407 => x"bd0bff88",
   408 => x"0c810ba0",
   409 => x"8093a858",
   410 => x"58835976",
   411 => x"08800c80",
   412 => x"08770856",
   413 => x"5473752e",
   414 => x"92388008",
   415 => x"537452a0",
   416 => x"8093b851",
   417 => x"a08080ed",
   418 => x"2d805880",
   419 => x"70575575",
   420 => x"70840557",
   421 => x"08811656",
   422 => x"54a08075",
   423 => x"24f13880",
   424 => x"08770856",
   425 => x"5675752e",
   426 => x"92388008",
   427 => x"537452a0",
   428 => x"8093f851",
   429 => x"a08080ed",
   430 => x"2d8058ff",
   431 => x"19841858",
   432 => x"59788025",
   433 => x"ffa53877",
   434 => x"802e8b38",
   435 => x"a08098b4",
   436 => x"51a08080",
   437 => x"ed2d8157",
   438 => x"85aad5aa",
   439 => x"d50b800c",
   440 => x"fad5aad5",
   441 => x"aa0b8c0c",
   442 => x"cc0b800b",
   443 => x"a08080b9",
   444 => x"2db30b8f",
   445 => x"0ba08080",
   446 => x"b92d8008",
   447 => x"5574fce2",
   448 => x"d5aad52e",
   449 => x"90388008",
   450 => x"52a08094",
   451 => x"b851a080",
   452 => x"80ed2d80",
   453 => x"578c0858",
   454 => x"77fad5aa",
   455 => x"d4b32e90",
   456 => x"388c0852",
   457 => x"a08094f4",
   458 => x"51a08080",
   459 => x"ed2d8057",
   460 => x"80705755",
   461 => x"75708405",
   462 => x"57088116",
   463 => x"5654a080",
   464 => x"7524f138",
   465 => x"80085978",
   466 => x"fce2d5aa",
   467 => x"d52e9038",
   468 => x"800852a0",
   469 => x"8095b051",
   470 => x"a08080ed",
   471 => x"2d80578c",
   472 => x"085473fa",
   473 => x"d5aad4b3",
   474 => x"2e80dd38",
   475 => x"8c0852a0",
   476 => x"8095ec51",
   477 => x"a08080ed",
   478 => x"2da08052",
   479 => x"8051a080",
   480 => x"8a832da0",
   481 => x"8099a408",
   482 => x"54a08099",
   483 => x"a408802e",
   484 => x"8b38a080",
   485 => x"98d851a0",
   486 => x"8080ed2d",
   487 => x"73528051",
   488 => x"a08087ed",
   489 => x"2da08099",
   490 => x"a408802e",
   491 => x"fdb338a0",
   492 => x"8098f051",
   493 => x"a08080ed",
   494 => x"2d810ba0",
   495 => x"8093a858",
   496 => x"588359a0",
   497 => x"808ceb04",
   498 => x"76802eff",
   499 => x"ac38a080",
   500 => x"998851a0",
   501 => x"8080ed2d",
   502 => x"a0808ef9",
   503 => x"04a08099",
   504 => x"b00802a0",
   505 => x"8099b00c",
   506 => x"fd3d0d80",
   507 => x"53a08099",
   508 => x"b0088c05",
   509 => x"0852a080",
   510 => x"99b00888",
   511 => x"05085180",
   512 => x"cf3fa080",
   513 => x"99a40870",
   514 => x"a08099a4",
   515 => x"0c54853d",
   516 => x"0da08099",
   517 => x"b00c04a0",
   518 => x"8099b008",
   519 => x"02a08099",
   520 => x"b00cfd3d",
   521 => x"0d8153a0",
   522 => x"8099b008",
   523 => x"8c050852",
   524 => x"a08099b0",
   525 => x"08880508",
   526 => x"51963fa0",
   527 => x"8099a408",
   528 => x"70a08099",
   529 => x"a40c5485",
   530 => x"3d0da080",
   531 => x"99b00c04",
   532 => x"a08099b0",
   533 => x"0802a080",
   534 => x"99b00cfd",
   535 => x"3d0d810b",
   536 => x"a08099b0",
   537 => x"08fc050c",
   538 => x"800ba080",
   539 => x"99b008f8",
   540 => x"050ca080",
   541 => x"99b0088c",
   542 => x"0508a080",
   543 => x"99b00888",
   544 => x"050827bf",
   545 => x"38a08099",
   546 => x"b008fc05",
   547 => x"08802eb3",
   548 => x"38800ba0",
   549 => x"8099b008",
   550 => x"8c050824",
   551 => x"a638a080",
   552 => x"99b0088c",
   553 => x"050810a0",
   554 => x"8099b008",
   555 => x"8c050ca0",
   556 => x"8099b008",
   557 => x"fc050810",
   558 => x"a08099b0",
   559 => x"08fc050c",
   560 => x"ffb039a0",
   561 => x"8099b008",
   562 => x"fc050880",
   563 => x"2e80ed38",
   564 => x"a08099b0",
   565 => x"088c0508",
   566 => x"a08099b0",
   567 => x"08880508",
   568 => x"26b338a0",
   569 => x"8099b008",
   570 => x"880508a0",
   571 => x"8099b008",
   572 => x"8c050831",
   573 => x"a08099b0",
   574 => x"0888050c",
   575 => x"a08099b0",
   576 => x"08f80508",
   577 => x"a08099b0",
   578 => x"08fc0508",
   579 => x"07a08099",
   580 => x"b008f805",
   581 => x"0ca08099",
   582 => x"b008fc05",
   583 => x"08812aa0",
   584 => x"8099b008",
   585 => x"fc050ca0",
   586 => x"8099b008",
   587 => x"8c050881",
   588 => x"2aa08099",
   589 => x"b0088c05",
   590 => x"0cff8839",
   591 => x"a08099b0",
   592 => x"08900508",
   593 => x"802e9538",
   594 => x"a08099b0",
   595 => x"08880508",
   596 => x"70a08099",
   597 => x"b008f405",
   598 => x"0c519339",
   599 => x"a08099b0",
   600 => x"08f80508",
   601 => x"70a08099",
   602 => x"b008f405",
   603 => x"0c51a080",
   604 => x"99b008f4",
   605 => x"0508a080",
   606 => x"99a40c85",
   607 => x"3d0da080",
   608 => x"99b00c04",
   609 => x"00ffffff",
   610 => x"ff00ffff",
   611 => x"ffff00ff",
   612 => x"ffffff00",
   613 => x"30313233",
   614 => x"34353637",
   615 => x"38394142",
   616 => x"43444546",
   617 => x"00000000",
   618 => x"00000000",
   619 => x"55555555",
   620 => x"aaaaaaaa",
   621 => x"ffffffff",
   622 => x"53616e69",
   623 => x"74792063",
   624 => x"6865636b",
   625 => x"20666169",
   626 => x"6c656420",
   627 => x"28626566",
   628 => x"6f726520",
   629 => x"63616368",
   630 => x"65207265",
   631 => x"66726573",
   632 => x"6829206f",
   633 => x"6e203078",
   634 => x"25642028",
   635 => x"676f7420",
   636 => x"30782564",
   637 => x"290a0000",
   638 => x"53616e69",
   639 => x"74792063",
   640 => x"6865636b",
   641 => x"20666169",
   642 => x"6c656420",
   643 => x"28616674",
   644 => x"65722063",
   645 => x"61636865",
   646 => x"20726566",
   647 => x"72657368",
   648 => x"29206f6e",
   649 => x"20307825",
   650 => x"64202867",
   651 => x"6f742030",
   652 => x"78256429",
   653 => x"0a000000",
   654 => x"42797465",
   655 => x"20636865",
   656 => x"636b2066",
   657 => x"61696c65",
   658 => x"64202862",
   659 => x"65666f72",
   660 => x"65206361",
   661 => x"63686520",
   662 => x"72656672",
   663 => x"65736829",
   664 => x"20617420",
   665 => x"30202867",
   666 => x"6f742030",
   667 => x"78256429",
   668 => x"0a000000",
   669 => x"42797465",
   670 => x"20636865",
   671 => x"636b2066",
   672 => x"61696c65",
   673 => x"64202862",
   674 => x"65666f72",
   675 => x"65206361",
   676 => x"63686520",
   677 => x"72656672",
   678 => x"65736829",
   679 => x"20617420",
   680 => x"33202867",
   681 => x"6f742030",
   682 => x"78256429",
   683 => x"0a000000",
   684 => x"42797465",
   685 => x"20636865",
   686 => x"636b2066",
   687 => x"61696c65",
   688 => x"64202861",
   689 => x"66746572",
   690 => x"20636163",
   691 => x"68652072",
   692 => x"65667265",
   693 => x"73682920",
   694 => x"61742030",
   695 => x"2028676f",
   696 => x"74203078",
   697 => x"2564290a",
   698 => x"00000000",
   699 => x"42797465",
   700 => x"20636865",
   701 => x"636b2066",
   702 => x"61696c65",
   703 => x"64202861",
   704 => x"66746572",
   705 => x"20636163",
   706 => x"68652072",
   707 => x"65667265",
   708 => x"73682920",
   709 => x"61742033",
   710 => x"2028676f",
   711 => x"74203078",
   712 => x"2564290a",
   713 => x"00000000",
   714 => x"43686563",
   715 => x"6b696e67",
   716 => x"206d656d",
   717 => x"6f727900",
   718 => x"30782564",
   719 => x"20676f6f",
   720 => x"64207265",
   721 => x"6164732c",
   722 => x"20000000",
   723 => x"4572726f",
   724 => x"72206174",
   725 => x"20307825",
   726 => x"642c2065",
   727 => x"78706563",
   728 => x"74656420",
   729 => x"30782564",
   730 => x"2c20676f",
   731 => x"74203078",
   732 => x"25640a00",
   733 => x"42616420",
   734 => x"64617461",
   735 => x"20666f75",
   736 => x"6e642061",
   737 => x"74203078",
   738 => x"25642028",
   739 => x"30782564",
   740 => x"290a0000",
   741 => x"53445241",
   742 => x"4d207369",
   743 => x"7a652028",
   744 => x"61737375",
   745 => x"6d696e67",
   746 => x"206e6f20",
   747 => x"61646472",
   748 => x"65737320",
   749 => x"6661756c",
   750 => x"74732920",
   751 => x"69732030",
   752 => x"78256420",
   753 => x"6d656761",
   754 => x"62797465",
   755 => x"730a0000",
   756 => x"416c6961",
   757 => x"73657320",
   758 => x"666f756e",
   759 => x"64206174",
   760 => x"20307825",
   761 => x"640a0000",
   762 => x"28416c69",
   763 => x"61736573",
   764 => x"2070726f",
   765 => x"6261626c",
   766 => x"79207369",
   767 => x"6d706c79",
   768 => x"20696e64",
   769 => x"69636174",
   770 => x"65207468",
   771 => x"61742052",
   772 => x"414d0a69",
   773 => x"7320736d",
   774 => x"616c6c65",
   775 => x"72207468",
   776 => x"616e2036",
   777 => x"34206d65",
   778 => x"67616279",
   779 => x"74657329",
   780 => x"0a000000",
   781 => x"46697273",
   782 => x"74207374",
   783 => x"61676520",
   784 => x"73616e69",
   785 => x"74792063",
   786 => x"6865636b",
   787 => x"20706173",
   788 => x"7365642e",
   789 => x"0a000000",
   790 => x"41646472",
   791 => x"65737320",
   792 => x"63686563",
   793 => x"6b207061",
   794 => x"73736564",
   795 => x"2e0a0000",
   796 => x"4c465352",
   797 => x"20636865",
   798 => x"636b2070",
   799 => x"61737365",
   800 => x"642e0a0a",
   801 => x"00000000",
   802 => x"42797465",
   803 => x"20286471",
   804 => x"6d292063",
   805 => x"6865636b",
   806 => x"20706173",
   807 => x"7365640a",
   808 => x"00000000",
	others => x"00000000"
);

begin

process (clk)
begin
	if (clk'event and clk = '1') then
		if (from_zpu.memAWriteEnable = '1') and (from_zpu.memBWriteEnable = '1') and (from_zpu.memAAddr=from_zpu.memBAddr) and (from_zpu.memAWrite/=from_zpu.memBWrite) then
			report "write collision" severity failure;
		end if;
	
		if (from_zpu.memAWriteEnable = '1') then
			ram(to_integer(unsigned(from_zpu.memAAddr(maxAddrBit downto 2)))) := from_zpu.memAWrite;
			to_zpu.memARead <= from_zpu.memAWrite;
		else
			to_zpu.memARead <= ram(to_integer(unsigned(from_zpu.memAAddr(maxAddrBit downto 2))));
		end if;
	end if;
end process;

process (clk)
begin
	if (clk'event and clk = '1') then
		if (from_zpu.memBWriteEnable = '1') then
			ram(to_integer(unsigned(from_zpu.memBAddr(maxAddrBit downto 2)))) := from_zpu.memBWrite;
			to_zpu.memBRead <= from_zpu.memBWrite;
		else
			to_zpu.memBRead <= ram(to_integer(unsigned(from_zpu.memBAddr(maxAddrBit downto 2))));
		end if;
	end if;
end process;


end arch;

