-- ZPU
--
-- Copyright 2004-2008 oharboe - �yvind Harboe - oyvind.harboe@zylin.com
-- Modified by Alastair M. Robinson for the ZPUFlex project.
--
-- The FreeBSD license
-- 
-- Redistribution and use in source and binary forms, with or without
-- modification, are permitted provided that the following conditions
-- are met:
-- 
-- 1. Redistributions of source code must retain the above copyright
--    notice, this list of conditions and the following disclaimer.
-- 2. Redistributions in binary form must reproduce the above
--    copyright notice, this list of conditions and the following
--    disclaimer in the documentation and/or other materials
--    provided with the distribution.
-- 
-- THIS SOFTWARE IS PROVIDED BY THE ZPU PROJECT ``AS IS'' AND ANY
-- EXPRESS OR IMPLIED WARRANTIES, INCLUDING, BUT NOT LIMITED TO,
-- THE IMPLIED WARRANTIES OF MERCHANTABILITY AND FITNESS FOR A
-- PARTICULAR PURPOSE ARE DISCLAIMED. IN NO EVENT SHALL THE
-- ZPU PROJECT OR CONTRIBUTORS BE LIABLE FOR ANY DIRECT,
-- INDIRECT, INCIDENTAL, SPECIAL, EXEMPLARY, OR CONSEQUENTIAL DAMAGES
-- (INCLUDING, BUT NOT LIMITED TO, PROCUREMENT OF SUBSTITUTE GOODS
-- OR SERVICES; LOSS OF USE, DATA, OR PROFITS; OR BUSINESS INTERRUPTION)
-- HOWEVER CAUSED AND ON ANY THEORY OF LIABILITY, WHETHER IN CONTRACT,
-- STRICT LIABILITY, OR TORT (INCLUDING NEGLIGENCE OR OTHERWISE)
-- ARISING IN ANY WAY OUT OF THE USE OF THIS SOFTWARE, EVEN IF
-- ADVISED OF THE POSSIBILITY OF SUCH DAMAGE.
-- 
-- The views and conclusions contained in the software and documentation
-- are those of the authors and should not be interpreted as representing
-- official policies, either expressed or implied, of the ZPU Project.

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;


library work;
use work.zpupkg.all;

entity Interrupt_ROM is
generic
	(
		maxAddrBitBRAM : integer := maxAddrBitBRAMLimit -- Specify your actual ROM size to save LEs and unnecessary block RAM usage.
	);
port (
	clk : in std_logic;
	areset : in std_logic := '0';
	from_zpu : in ZPU_ToROM;
	to_zpu : out ZPU_FromROM
);
end Interrupt_ROM;

architecture arch of Interrupt_ROM is

type ram_type is array(natural range 0 to ((2**(maxAddrBitBRAM+1))/4)-1) of std_logic_vector(wordSize-1 downto 0);

shared variable ram : ram_type :=
(
     0 => x"0b0b0b88",
     1 => x"e5040000",
     2 => x"00000000",
     3 => x"00000000",
     4 => x"00000000",
     5 => x"00000000",
     6 => x"00000000",
     7 => x"00000000",
     8 => x"88088c08",
     9 => x"90080b0b",
    10 => x"0b88e108",
    11 => x"2d900c8c",
    12 => x"0c880c04",
    13 => x"00000000",
    14 => x"00000000",
    15 => x"00000000",
    16 => x"71fd0608",
    17 => x"72830609",
    18 => x"81058205",
    19 => x"832b2a83",
    20 => x"ffff0652",
    21 => x"04000000",
    22 => x"00000000",
    23 => x"00000000",
    24 => x"71fd0608",
    25 => x"83ffff73",
    26 => x"83060981",
    27 => x"05820583",
    28 => x"2b2b0906",
    29 => x"7383ffff",
    30 => x"0b0b0b0b",
    31 => x"83a50400",
    32 => x"72098105",
    33 => x"72057373",
    34 => x"09060906",
    35 => x"73097306",
    36 => x"070a8106",
    37 => x"53510400",
    38 => x"00000000",
    39 => x"00000000",
    40 => x"72722473",
    41 => x"732e0753",
    42 => x"51040000",
    43 => x"00000000",
    44 => x"00000000",
    45 => x"00000000",
    46 => x"00000000",
    47 => x"00000000",
    48 => x"71737109",
    49 => x"71068106",
    50 => x"09810572",
    51 => x"0a100a72",
    52 => x"0a100a31",
    53 => x"050a8106",
    54 => x"51515351",
    55 => x"04000000",
    56 => x"72722673",
    57 => x"732e0753",
    58 => x"51040000",
    59 => x"00000000",
    60 => x"00000000",
    61 => x"00000000",
    62 => x"00000000",
    63 => x"00000000",
    64 => x"00000000",
    65 => x"00000000",
    66 => x"00000000",
    67 => x"00000000",
    68 => x"00000000",
    69 => x"00000000",
    70 => x"00000000",
    71 => x"00000000",
    72 => x"0b0b0b88",
    73 => x"ba040000",
    74 => x"00000000",
    75 => x"00000000",
    76 => x"00000000",
    77 => x"00000000",
    78 => x"00000000",
    79 => x"00000000",
    80 => x"720a722b",
    81 => x"0a535104",
    82 => x"00000000",
    83 => x"00000000",
    84 => x"00000000",
    85 => x"00000000",
    86 => x"00000000",
    87 => x"00000000",
    88 => x"72729f06",
    89 => x"0981050b",
    90 => x"0b0b889f",
    91 => x"05040000",
    92 => x"00000000",
    93 => x"00000000",
    94 => x"00000000",
    95 => x"00000000",
    96 => x"72722aff",
    97 => x"739f062a",
    98 => x"0974090a",
    99 => x"8106ff05",
   100 => x"06075351",
   101 => x"04000000",
   102 => x"00000000",
   103 => x"00000000",
   104 => x"71715351",
   105 => x"04067383",
   106 => x"06098105",
   107 => x"8205832b",
   108 => x"0b2b0772",
   109 => x"fc060c51",
   110 => x"51040000",
   111 => x"00000000",
   112 => x"72098105",
   113 => x"72050970",
   114 => x"81050906",
   115 => x"0a810653",
   116 => x"51040000",
   117 => x"00000000",
   118 => x"00000000",
   119 => x"00000000",
   120 => x"72098105",
   121 => x"72050970",
   122 => x"81050906",
   123 => x"0a098106",
   124 => x"53510400",
   125 => x"00000000",
   126 => x"00000000",
   127 => x"00000000",
   128 => x"71098105",
   129 => x"52040000",
   130 => x"00000000",
   131 => x"00000000",
   132 => x"00000000",
   133 => x"00000000",
   134 => x"00000000",
   135 => x"00000000",
   136 => x"72720981",
   137 => x"05055351",
   138 => x"04000000",
   139 => x"00000000",
   140 => x"00000000",
   141 => x"00000000",
   142 => x"00000000",
   143 => x"00000000",
   144 => x"72097206",
   145 => x"73730906",
   146 => x"07535104",
   147 => x"00000000",
   148 => x"00000000",
   149 => x"00000000",
   150 => x"00000000",
   151 => x"00000000",
   152 => x"71fc0608",
   153 => x"72830609",
   154 => x"81058305",
   155 => x"1010102a",
   156 => x"81ff0652",
   157 => x"04000000",
   158 => x"00000000",
   159 => x"00000000",
   160 => x"71fc0608",
   161 => x"0b0b0b91",
   162 => x"b0738306",
   163 => x"10100508",
   164 => x"060b0b0b",
   165 => x"88a20400",
   166 => x"00000000",
   167 => x"00000000",
   168 => x"88088c08",
   169 => x"90087575",
   170 => x"0b0b0b8d",
   171 => x"b12d5050",
   172 => x"88085690",
   173 => x"0c8c0c88",
   174 => x"0c510400",
   175 => x"00000000",
   176 => x"88088c08",
   177 => x"90087575",
   178 => x"0b0b0b8e",
   179 => x"e32d5050",
   180 => x"88085690",
   181 => x"0c8c0c88",
   182 => x"0c510400",
   183 => x"00000000",
   184 => x"72097081",
   185 => x"0509060a",
   186 => x"8106ff05",
   187 => x"70547106",
   188 => x"73097274",
   189 => x"05ff0506",
   190 => x"07515151",
   191 => x"04000000",
   192 => x"72097081",
   193 => x"0509060a",
   194 => x"098106ff",
   195 => x"05705471",
   196 => x"06730972",
   197 => x"7405ff05",
   198 => x"06075151",
   199 => x"51040000",
   200 => x"05ff0504",
   201 => x"00000000",
   202 => x"00000000",
   203 => x"00000000",
   204 => x"00000000",
   205 => x"00000000",
   206 => x"00000000",
   207 => x"00000000",
   208 => x"04000000",
   209 => x"00000000",
   210 => x"00000000",
   211 => x"00000000",
   212 => x"00000000",
   213 => x"00000000",
   214 => x"00000000",
   215 => x"00000000",
   216 => x"71810552",
   217 => x"04000000",
   218 => x"00000000",
   219 => x"00000000",
   220 => x"00000000",
   221 => x"00000000",
   222 => x"00000000",
   223 => x"00000000",
   224 => x"04000000",
   225 => x"00000000",
   226 => x"00000000",
   227 => x"00000000",
   228 => x"00000000",
   229 => x"00000000",
   230 => x"00000000",
   231 => x"00000000",
   232 => x"02840572",
   233 => x"10100552",
   234 => x"04000000",
   235 => x"00000000",
   236 => x"00000000",
   237 => x"00000000",
   238 => x"00000000",
   239 => x"00000000",
   240 => x"00000000",
   241 => x"00000000",
   242 => x"00000000",
   243 => x"00000000",
   244 => x"00000000",
   245 => x"00000000",
   246 => x"00000000",
   247 => x"00000000",
   248 => x"717105ff",
   249 => x"05715351",
   250 => x"020d0400",
   251 => x"00000000",
   252 => x"00000000",
   253 => x"00000000",
   254 => x"00000000",
   255 => x"00000000",
   256 => x"10101010",
   257 => x"10101010",
   258 => x"10101010",
   259 => x"10101010",
   260 => x"10101010",
   261 => x"10101010",
   262 => x"10101010",
   263 => x"10101053",
   264 => x"51047381",
   265 => x"ff067383",
   266 => x"06098105",
   267 => x"83051010",
   268 => x"102b0772",
   269 => x"fc060c51",
   270 => x"51047272",
   271 => x"80728106",
   272 => x"ff050972",
   273 => x"06057110",
   274 => x"52720a10",
   275 => x"0a5372ed",
   276 => x"38515153",
   277 => x"51040000",
   278 => x"80040088",
   279 => x"da040400",
   280 => x"00000004",
   281 => x"5e92b070",
   282 => x"93c4278b",
   283 => x"38807170",
   284 => x"8405530c",
   285 => x"88e70488",
   286 => x"da518cfb",
   287 => x"04f93d0d",
   288 => x"797b7d0b",
   289 => x"0b0b92b0",
   290 => x"585a5754",
   291 => x"80577377",
   292 => x"258938ad",
   293 => x"5182c23f",
   294 => x"73305473",
   295 => x"8e38b00b",
   296 => x"0b0b0b92",
   297 => x"b0348115",
   298 => x"55a03977",
   299 => x"743691c0",
   300 => x"05537233",
   301 => x"75708105",
   302 => x"57347774",
   303 => x"355473eb",
   304 => x"38740b0b",
   305 => x"0b92b02e",
   306 => x"9138ff15",
   307 => x"55743376",
   308 => x"70810558",
   309 => x"34811757",
   310 => x"e8398076",
   311 => x"3476880c",
   312 => x"893d0d04",
   313 => x"f13d0d92",
   314 => x"3d578070",
   315 => x"78708405",
   316 => x"5a087241",
   317 => x"5f5d587c",
   318 => x"7084055e",
   319 => x"085a805b",
   320 => x"79982a7a",
   321 => x"882b5b56",
   322 => x"75863877",
   323 => x"5f81c339",
   324 => x"7d802e81",
   325 => x"9d38805e",
   326 => x"7580e42e",
   327 => x"8a387580",
   328 => x"f82e0981",
   329 => x"06893876",
   330 => x"84187108",
   331 => x"5e585475",
   332 => x"80e42e9e",
   333 => x"387580e4",
   334 => x"268a3875",
   335 => x"80e32ebf",
   336 => x"3880c639",
   337 => x"7580f32e",
   338 => x"a5387580",
   339 => x"f82e8738",
   340 => x"b8398a53",
   341 => x"83399053",
   342 => x"0b0b0b93",
   343 => x"80527b51",
   344 => x"fe9b3f88",
   345 => x"080b0b0b",
   346 => x"93805a55",
   347 => x"ab397684",
   348 => x"18710870",
   349 => x"545b5854",
   350 => x"80fe3f80",
   351 => x"559a3976",
   352 => x"84187108",
   353 => x"585854b6",
   354 => x"39a55180",
   355 => x"cc3f7551",
   356 => x"80c73f82",
   357 => x"1858ae39",
   358 => x"74ff1656",
   359 => x"54807425",
   360 => x"a4387870",
   361 => x"81055a33",
   362 => x"705256ad",
   363 => x"3f811858",
   364 => x"e73975a5",
   365 => x"2e098106",
   366 => x"8538815e",
   367 => x"88397551",
   368 => x"983f8118",
   369 => x"58811b5b",
   370 => x"837b25fe",
   371 => x"b33875fe",
   372 => x"a6387e88",
   373 => x"0c913d0d",
   374 => x"04ff3d0d",
   375 => x"7352c008",
   376 => x"70882a70",
   377 => x"81065151",
   378 => x"5170802e",
   379 => x"f13871c0",
   380 => x"0c71880c",
   381 => x"833d0d04",
   382 => x"fb3d0d80",
   383 => x"78575575",
   384 => x"70840557",
   385 => x"08538054",
   386 => x"72982a73",
   387 => x"882b5452",
   388 => x"71802ea2",
   389 => x"38c00870",
   390 => x"882a7081",
   391 => x"06515151",
   392 => x"70802ef1",
   393 => x"3871c00c",
   394 => x"81158115",
   395 => x"55558374",
   396 => x"25d63871",
   397 => x"ca387488",
   398 => x"0c873d0d",
   399 => x"047188e1",
   400 => x"0c04ffb0",
   401 => x"08880c04",
   402 => x"810bffb0",
   403 => x"0c04800b",
   404 => x"ffb00c04",
   405 => x"ff3d0df6",
   406 => x"3fe83f93",
   407 => x"c0088132",
   408 => x"7093c00c",
   409 => x"5271802e",
   410 => x"863891d4",
   411 => x"51843991",
   412 => x"e051ff84",
   413 => x"3fd23f83",
   414 => x"3d0d0480",
   415 => x"3d0d800b",
   416 => x"93c00c91",
   417 => x"ec51fef0",
   418 => x"3f800bf8",
   419 => x"840c868d",
   420 => x"a00bf888",
   421 => x"0c928451",
   422 => x"fede3f8c",
   423 => x"d451ff9d",
   424 => x"3fffa53f",
   425 => x"929c51fe",
   426 => x"cf3f810b",
   427 => x"f8800cff",
   428 => x"39940802",
   429 => x"940cf93d",
   430 => x"0d800b94",
   431 => x"08fc050c",
   432 => x"94088805",
   433 => x"088025ab",
   434 => x"38940888",
   435 => x"05083094",
   436 => x"0888050c",
   437 => x"800b9408",
   438 => x"f4050c94",
   439 => x"08fc0508",
   440 => x"8838810b",
   441 => x"9408f405",
   442 => x"0c9408f4",
   443 => x"05089408",
   444 => x"fc050c94",
   445 => x"088c0508",
   446 => x"8025ab38",
   447 => x"94088c05",
   448 => x"08309408",
   449 => x"8c050c80",
   450 => x"0b9408f0",
   451 => x"050c9408",
   452 => x"fc050888",
   453 => x"38810b94",
   454 => x"08f0050c",
   455 => x"9408f005",
   456 => x"089408fc",
   457 => x"050c8053",
   458 => x"94088c05",
   459 => x"08529408",
   460 => x"88050851",
   461 => x"81a73f88",
   462 => x"08709408",
   463 => x"f8050c54",
   464 => x"9408fc05",
   465 => x"08802e8c",
   466 => x"389408f8",
   467 => x"05083094",
   468 => x"08f8050c",
   469 => x"9408f805",
   470 => x"0870880c",
   471 => x"54893d0d",
   472 => x"940c0494",
   473 => x"0802940c",
   474 => x"fb3d0d80",
   475 => x"0b9408fc",
   476 => x"050c9408",
   477 => x"88050880",
   478 => x"25933894",
   479 => x"08880508",
   480 => x"30940888",
   481 => x"050c810b",
   482 => x"9408fc05",
   483 => x"0c94088c",
   484 => x"05088025",
   485 => x"8c389408",
   486 => x"8c050830",
   487 => x"94088c05",
   488 => x"0c815394",
   489 => x"088c0508",
   490 => x"52940888",
   491 => x"050851ad",
   492 => x"3f880870",
   493 => x"9408f805",
   494 => x"0c549408",
   495 => x"fc050880",
   496 => x"2e8c3894",
   497 => x"08f80508",
   498 => x"309408f8",
   499 => x"050c9408",
   500 => x"f8050870",
   501 => x"880c5487",
   502 => x"3d0d940c",
   503 => x"04940802",
   504 => x"940cfd3d",
   505 => x"0d810b94",
   506 => x"08fc050c",
   507 => x"800b9408",
   508 => x"f8050c94",
   509 => x"088c0508",
   510 => x"94088805",
   511 => x"0827ac38",
   512 => x"9408fc05",
   513 => x"08802ea3",
   514 => x"38800b94",
   515 => x"088c0508",
   516 => x"24993894",
   517 => x"088c0508",
   518 => x"1094088c",
   519 => x"050c9408",
   520 => x"fc050810",
   521 => x"9408fc05",
   522 => x"0cc93994",
   523 => x"08fc0508",
   524 => x"802e80c9",
   525 => x"3894088c",
   526 => x"05089408",
   527 => x"88050826",
   528 => x"a1389408",
   529 => x"88050894",
   530 => x"088c0508",
   531 => x"31940888",
   532 => x"050c9408",
   533 => x"f8050894",
   534 => x"08fc0508",
   535 => x"079408f8",
   536 => x"050c9408",
   537 => x"fc050881",
   538 => x"2a9408fc",
   539 => x"050c9408",
   540 => x"8c050881",
   541 => x"2a94088c",
   542 => x"050cffaf",
   543 => x"39940890",
   544 => x"0508802e",
   545 => x"8f389408",
   546 => x"88050870",
   547 => x"9408f405",
   548 => x"0c518d39",
   549 => x"9408f805",
   550 => x"08709408",
   551 => x"f4050c51",
   552 => x"9408f405",
   553 => x"08880c85",
   554 => x"3d0d940c",
   555 => x"04000000",
   556 => x"00ffffff",
   557 => x"ff00ffff",
   558 => x"ffff00ff",
   559 => x"ffffff00",
   560 => x"30313233",
   561 => x"34353637",
   562 => x"38394142",
   563 => x"43444546",
   564 => x"00000000",
   565 => x"5469636b",
   566 => x"2e2e2e0a",
   567 => x"00000000",
   568 => x"546f636b",
   569 => x"2e2e2e0a",
   570 => x"00000000",
   571 => x"53657474",
   572 => x"696e6720",
   573 => x"75702074",
   574 => x"696d6572",
   575 => x"2e2e2e0a",
   576 => x"00000000",
   577 => x"456e6162",
   578 => x"6c696e67",
   579 => x"20696e74",
   580 => x"65727275",
   581 => x"7074732e",
   582 => x"2e2e0a00",
   583 => x"456e6162",
   584 => x"6c696e67",
   585 => x"2074696d",
   586 => x"65722e2e",
   587 => x"2e0a002e",
	others => x"00000000"
);

begin

process (clk)
begin
	if (clk'event and clk = '1') then
		if (from_zpu.memAWriteEnable = '1') and (from_zpu.memBWriteEnable = '1') and (from_zpu.memAAddr=from_zpu.memBAddr) and (from_zpu.memAWrite/=from_zpu.memBWrite) then
			report "write collision" severity failure;
		end if;
	
		if (from_zpu.memAWriteEnable = '1') then
			ram(to_integer(unsigned(from_zpu.memAAddr(maxAddrBitBRAM downto 2)))) := from_zpu.memAWrite;
			to_zpu.memARead <= from_zpu.memAWrite;
		else
			to_zpu.memARead <= ram(to_integer(unsigned(from_zpu.memAAddr(maxAddrBitBRAM downto 2))));
		end if;
	end if;
end process;

process (clk)
begin
	if (clk'event and clk = '1') then
		if (from_zpu.memBWriteEnable = '1') then
			ram(to_integer(unsigned(from_zpu.memBAddr(maxAddrBitBRAM downto 2)))) := from_zpu.memBWrite;
			to_zpu.memBRead <= from_zpu.memBWrite;
		else
			to_zpu.memBRead <= ram(to_integer(unsigned(from_zpu.memBAddr(maxAddrBitBRAM downto 2))));
		end if;
	end if;
end process;


end arch;

