-- ZPU
--
-- Copyright 2004-2008 oharboe - �yvind Harboe - oyvind.harboe@zylin.com
-- Modified by Alastair M. Robinson for the ZPUFlex project.
--
-- The FreeBSD license
-- 
-- Redistribution and use in source and binary forms, with or without
-- modification, are permitted provided that the following conditions
-- are met:
-- 
-- 1. Redistributions of source code must retain the above copyright
--    notice, this list of conditions and the following disclaimer.
-- 2. Redistributions in binary form must reproduce the above
--    copyright notice, this list of conditions and the following
--    disclaimer in the documentation and/or other materials
--    provided with the distribution.
-- 
-- THIS SOFTWARE IS PROVIDED BY THE ZPU PROJECT ``AS IS'' AND ANY
-- EXPRESS OR IMPLIED WARRANTIES, INCLUDING, BUT NOT LIMITED TO,
-- THE IMPLIED WARRANTIES OF MERCHANTABILITY AND FITNESS FOR A
-- PARTICULAR PURPOSE ARE DISCLAIMED. IN NO EVENT SHALL THE
-- ZPU PROJECT OR CONTRIBUTORS BE LIABLE FOR ANY DIRECT,
-- INDIRECT, INCIDENTAL, SPECIAL, EXEMPLARY, OR CONSEQUENTIAL DAMAGES
-- (INCLUDING, BUT NOT LIMITED TO, PROCUREMENT OF SUBSTITUTE GOODS
-- OR SERVICES; LOSS OF USE, DATA, OR PROFITS; OR BUSINESS INTERRUPTION)
-- HOWEVER CAUSED AND ON ANY THEORY OF LIABILITY, WHETHER IN CONTRACT,
-- STRICT LIABILITY, OR TORT (INCLUDING NEGLIGENCE OR OTHERWISE)
-- ARISING IN ANY WAY OUT OF THE USE OF THIS SOFTWARE, EVEN IF
-- ADVISED OF THE POSSIBILITY OF SUCH DAMAGE.
-- 
-- The views and conclusions contained in the software and documentation
-- are those of the authors and should not be interpreted as representing
-- official policies, either expressed or implied, of the ZPU Project.

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;


library work;
use work.zpu_config.all;
use work.zpupkg.all;

entity Dhrystone_min_ROM is
generic
	(
		maxAddrBitBRAM : integer := maxAddrBitBRAMLimit -- Specify your actual ROM size to save LEs and unnecessary block RAM usage.
	);
port (
	clk : in std_logic;
	areset : in std_logic := '0';
	from_zpu : in ZPU_ToROM;
	to_zpu : out ZPU_FromROM
);
end Dhrystone_min_ROM;

architecture arch of Dhrystone_min_ROM is

type ram_type is array(natural range 0 to ((2**(maxAddrBitBRAM+1))/4)-1) of std_logic_vector(wordSize-1 downto 0);

shared variable ram : ram_type :=
(
     0 => x"0b0b0b88",
     1 => x"dd040000",
     2 => x"00000000",
     3 => x"00000000",
     4 => x"00000000",
     5 => x"00000000",
     6 => x"00000000",
     7 => x"00000000",
     8 => x"88088c08",
     9 => x"90080b0b",
    10 => x"0b88e708",
    11 => x"2d900c8c",
    12 => x"0c880c04",
    13 => x"00000000",
    14 => x"00000000",
    15 => x"00000000",
    16 => x"71fd0608",
    17 => x"72830609",
    18 => x"81058205",
    19 => x"832b2a83",
    20 => x"ffff0652",
    21 => x"04000000",
    22 => x"00000000",
    23 => x"00000000",
    24 => x"71fd0608",
    25 => x"83ffff73",
    26 => x"83060981",
    27 => x"05820583",
    28 => x"2b2b0906",
    29 => x"7383ffff",
    30 => x"0b0b0b0b",
    31 => x"83a50400",
    32 => x"72098105",
    33 => x"72057373",
    34 => x"09060906",
    35 => x"73097306",
    36 => x"070a8106",
    37 => x"53510400",
    38 => x"00000000",
    39 => x"00000000",
    40 => x"72722473",
    41 => x"732e0753",
    42 => x"51040000",
    43 => x"00000000",
    44 => x"00000000",
    45 => x"00000000",
    46 => x"00000000",
    47 => x"00000000",
    48 => x"71737109",
    49 => x"71068106",
    50 => x"09810572",
    51 => x"0a100a72",
    52 => x"0a100a31",
    53 => x"050a8106",
    54 => x"51515351",
    55 => x"04000000",
    56 => x"72722673",
    57 => x"732e0753",
    58 => x"51040000",
    59 => x"00000000",
    60 => x"00000000",
    61 => x"00000000",
    62 => x"00000000",
    63 => x"00000000",
    64 => x"00000000",
    65 => x"00000000",
    66 => x"00000000",
    67 => x"00000000",
    68 => x"00000000",
    69 => x"00000000",
    70 => x"00000000",
    71 => x"00000000",
    72 => x"0b0b0b88",
    73 => x"ba040000",
    74 => x"00000000",
    75 => x"00000000",
    76 => x"00000000",
    77 => x"00000000",
    78 => x"00000000",
    79 => x"00000000",
    80 => x"720a722b",
    81 => x"0a535104",
    82 => x"00000000",
    83 => x"00000000",
    84 => x"00000000",
    85 => x"00000000",
    86 => x"00000000",
    87 => x"00000000",
    88 => x"72729f06",
    89 => x"0981050b",
    90 => x"0b0b889f",
    91 => x"05040000",
    92 => x"00000000",
    93 => x"00000000",
    94 => x"00000000",
    95 => x"00000000",
    96 => x"72722aff",
    97 => x"739f062a",
    98 => x"0974090a",
    99 => x"8106ff05",
   100 => x"06075351",
   101 => x"04000000",
   102 => x"00000000",
   103 => x"00000000",
   104 => x"71715351",
   105 => x"04067383",
   106 => x"06098105",
   107 => x"8205832b",
   108 => x"0b2b0772",
   109 => x"fc060c51",
   110 => x"51040000",
   111 => x"00000000",
   112 => x"72098105",
   113 => x"72050970",
   114 => x"81050906",
   115 => x"0a810653",
   116 => x"51040000",
   117 => x"00000000",
   118 => x"00000000",
   119 => x"00000000",
   120 => x"72098105",
   121 => x"72050970",
   122 => x"81050906",
   123 => x"0a098106",
   124 => x"53510400",
   125 => x"00000000",
   126 => x"00000000",
   127 => x"00000000",
   128 => x"71098105",
   129 => x"52040000",
   130 => x"00000000",
   131 => x"00000000",
   132 => x"00000000",
   133 => x"00000000",
   134 => x"00000000",
   135 => x"00000000",
   136 => x"72720981",
   137 => x"05055351",
   138 => x"04000000",
   139 => x"00000000",
   140 => x"00000000",
   141 => x"00000000",
   142 => x"00000000",
   143 => x"00000000",
   144 => x"72097206",
   145 => x"73730906",
   146 => x"07535104",
   147 => x"00000000",
   148 => x"00000000",
   149 => x"00000000",
   150 => x"00000000",
   151 => x"00000000",
   152 => x"71fc0608",
   153 => x"72830609",
   154 => x"81058305",
   155 => x"1010102a",
   156 => x"81ff0652",
   157 => x"04000000",
   158 => x"00000000",
   159 => x"00000000",
   160 => x"71fc0608",
   161 => x"0b0b0ba0",
   162 => x"84738306",
   163 => x"10100508",
   164 => x"060b0b0b",
   165 => x"88a20400",
   166 => x"00000000",
   167 => x"00000000",
   168 => x"88088c08",
   169 => x"90087575",
   170 => x"0b0b0b98",
   171 => x"f82d5050",
   172 => x"88085690",
   173 => x"0c8c0c88",
   174 => x"0c510400",
   175 => x"00000000",
   176 => x"88088c08",
   177 => x"90087575",
   178 => x"0b0b0b9a",
   179 => x"aa2d5050",
   180 => x"88085690",
   181 => x"0c8c0c88",
   182 => x"0c510400",
   183 => x"00000000",
   184 => x"72097081",
   185 => x"0509060a",
   186 => x"8106ff05",
   187 => x"70547106",
   188 => x"73097274",
   189 => x"05ff0506",
   190 => x"07515151",
   191 => x"04000000",
   192 => x"72097081",
   193 => x"0509060a",
   194 => x"098106ff",
   195 => x"05705471",
   196 => x"06730972",
   197 => x"7405ff05",
   198 => x"06075151",
   199 => x"51040000",
   200 => x"05ff0504",
   201 => x"00000000",
   202 => x"00000000",
   203 => x"00000000",
   204 => x"00000000",
   205 => x"00000000",
   206 => x"00000000",
   207 => x"00000000",
   208 => x"04000000",
   209 => x"00000000",
   210 => x"00000000",
   211 => x"00000000",
   212 => x"00000000",
   213 => x"00000000",
   214 => x"00000000",
   215 => x"00000000",
   216 => x"71810552",
   217 => x"04000000",
   218 => x"00000000",
   219 => x"00000000",
   220 => x"00000000",
   221 => x"00000000",
   222 => x"00000000",
   223 => x"00000000",
   224 => x"00000000",
   225 => x"00000000",
   226 => x"00000000",
   227 => x"00000000",
   228 => x"00000000",
   229 => x"00000000",
   230 => x"00000000",
   231 => x"00000000",
   232 => x"02840572",
   233 => x"10100552",
   234 => x"04000000",
   235 => x"00000000",
   236 => x"00000000",
   237 => x"00000000",
   238 => x"00000000",
   239 => x"00000000",
   240 => x"00000000",
   241 => x"00000000",
   242 => x"00000000",
   243 => x"00000000",
   244 => x"00000000",
   245 => x"00000000",
   246 => x"00000000",
   247 => x"00000000",
   248 => x"717105ff",
   249 => x"05715351",
   250 => x"020d0400",
   251 => x"00000000",
   252 => x"00000000",
   253 => x"00000000",
   254 => x"00000000",
   255 => x"00000000",
   256 => x"10101010",
   257 => x"10101010",
   258 => x"10101010",
   259 => x"10101010",
   260 => x"10101010",
   261 => x"10101010",
   262 => x"10101010",
   263 => x"10101053",
   264 => x"51047381",
   265 => x"ff067383",
   266 => x"06098105",
   267 => x"83051010",
   268 => x"102b0772",
   269 => x"fc060c51",
   270 => x"51047272",
   271 => x"80728106",
   272 => x"ff050972",
   273 => x"06057110",
   274 => x"52720a10",
   275 => x"0a5372ed",
   276 => x"38515153",
   277 => x"51040000",
   278 => x"800488da",
   279 => x"0488da0b",
   280 => x"8f820404",
   281 => x"00000000",
   282 => x"000463f1",
   283 => x"3d0d923d",
   284 => x"0b0b0ba5",
   285 => x"ac5a5c80",
   286 => x"7c708405",
   287 => x"5e08715f",
   288 => x"5f577d70",
   289 => x"84055f08",
   290 => x"56805875",
   291 => x"982a7688",
   292 => x"2b575574",
   293 => x"802e82b5",
   294 => x"387c802e",
   295 => x"b738805d",
   296 => x"7480e42e",
   297 => x"81983874",
   298 => x"80e42680",
   299 => x"d8387480",
   300 => x"e32eb738",
   301 => x"a551829c",
   302 => x"3f745182",
   303 => x"973f8217",
   304 => x"57811858",
   305 => x"837825c3",
   306 => x"3874ffb6",
   307 => x"387e880c",
   308 => x"913d0d04",
   309 => x"74a52e09",
   310 => x"81069738",
   311 => x"810b8119",
   312 => x"595d8378",
   313 => x"25ffa438",
   314 => x"e0397b84",
   315 => x"1d710857",
   316 => x"5d5a7451",
   317 => x"81de3f81",
   318 => x"17811959",
   319 => x"57837825",
   320 => x"ff8938c5",
   321 => x"397480f3",
   322 => x"2e098106",
   323 => x"ffa6387b",
   324 => x"841d7108",
   325 => x"70545b5d",
   326 => x"5481d83f",
   327 => x"800bff11",
   328 => x"55538073",
   329 => x"25ff9a38",
   330 => x"78708105",
   331 => x"5a337052",
   332 => x"5581a13f",
   333 => x"811774ff",
   334 => x"16565457",
   335 => x"e5397b84",
   336 => x"1d71080b",
   337 => x"0b0ba5ac",
   338 => x"0b0b0b0b",
   339 => x"a4dc615f",
   340 => x"585e525d",
   341 => x"5372b138",
   342 => x"b00b0b0b",
   343 => x"0ba4dc34",
   344 => x"811454ff",
   345 => x"14547333",
   346 => x"7b708105",
   347 => x"5d34811a",
   348 => x"5a730b0b",
   349 => x"0ba4dc2e",
   350 => x"098106e7",
   351 => x"38807b34",
   352 => x"79ff1155",
   353 => x"53ff9b39",
   354 => x"8a527251",
   355 => x"8dc53f88",
   356 => x"08a09405",
   357 => x"33747081",
   358 => x"0556348a",
   359 => x"5272518d",
   360 => x"8d3f8808",
   361 => x"538808e0",
   362 => x"38730b0b",
   363 => x"0ba4dc2e",
   364 => x"cc38ff14",
   365 => x"5473337b",
   366 => x"7081055d",
   367 => x"34811a5a",
   368 => x"730b0b0b",
   369 => x"a4dc2eff",
   370 => x"b438ff97",
   371 => x"3976880c",
   372 => x"913d0d04",
   373 => x"ff3d0d73",
   374 => x"52c00870",
   375 => x"882a7081",
   376 => x"06515151",
   377 => x"70802ef1",
   378 => x"3871c00c",
   379 => x"71880c83",
   380 => x"3d0d04fb",
   381 => x"3d0d8078",
   382 => x"57557570",
   383 => x"84055708",
   384 => x"53805472",
   385 => x"982a7388",
   386 => x"2b545271",
   387 => x"802ea238",
   388 => x"c0087088",
   389 => x"2a708106",
   390 => x"51515170",
   391 => x"802ef138",
   392 => x"71c00c81",
   393 => x"15811555",
   394 => x"55837425",
   395 => x"d63871ca",
   396 => x"3874880c",
   397 => x"873d0d04",
   398 => x"803d0dc8",
   399 => x"08f88011",
   400 => x"08880c51",
   401 => x"823d0d04",
   402 => x"803d0d80",
   403 => x"c10b80f4",
   404 => x"f834800b",
   405 => x"80f7900c",
   406 => x"70880c82",
   407 => x"3d0d04ff",
   408 => x"3d0d800b",
   409 => x"80f4f833",
   410 => x"52527080",
   411 => x"c12e9938",
   412 => x"7180f790",
   413 => x"080780f7",
   414 => x"900c80c2",
   415 => x"0b80f4fc",
   416 => x"3470880c",
   417 => x"833d0d04",
   418 => x"810b80f7",
   419 => x"90080780",
   420 => x"f7900c80",
   421 => x"c20b80f4",
   422 => x"fc347088",
   423 => x"0c833d0d",
   424 => x"04fd3d0d",
   425 => x"7570088a",
   426 => x"05535380",
   427 => x"f4f83351",
   428 => x"7080c12e",
   429 => x"8b3873f3",
   430 => x"3870880c",
   431 => x"853d0d04",
   432 => x"ff127080",
   433 => x"f4f40831",
   434 => x"740c880c",
   435 => x"853d0d04",
   436 => x"fc3d0d80",
   437 => x"f5a00855",
   438 => x"74802e8c",
   439 => x"38767508",
   440 => x"710c80f5",
   441 => x"a0085654",
   442 => x"8c155380",
   443 => x"f4f40852",
   444 => x"8a5188a7",
   445 => x"3f73880c",
   446 => x"863d0d04",
   447 => x"fb3d0d77",
   448 => x"70085656",
   449 => x"b05380f5",
   450 => x"a0085274",
   451 => x"518fc73f",
   452 => x"850b8c17",
   453 => x"0c850b8c",
   454 => x"160c7508",
   455 => x"750c80f5",
   456 => x"a0085473",
   457 => x"802e8a38",
   458 => x"7308750c",
   459 => x"80f5a008",
   460 => x"548c1453",
   461 => x"80f4f408",
   462 => x"528a5187",
   463 => x"de3f8415",
   464 => x"08ad3886",
   465 => x"0b8c160c",
   466 => x"88155288",
   467 => x"16085186",
   468 => x"ea3f80f5",
   469 => x"a0087008",
   470 => x"760c548c",
   471 => x"15705454",
   472 => x"8a527308",
   473 => x"5187b43f",
   474 => x"73880c87",
   475 => x"3d0d0475",
   476 => x"0854b053",
   477 => x"73527551",
   478 => x"8edc3f73",
   479 => x"880c873d",
   480 => x"0d04f33d",
   481 => x"0d80f48c",
   482 => x"0b80f4c0",
   483 => x"0c80f4c4",
   484 => x"0b80f5a0",
   485 => x"0c80f48c",
   486 => x"0b80f4c4",
   487 => x"0c800b80",
   488 => x"f4c40b84",
   489 => x"050c820b",
   490 => x"80f4c40b",
   491 => x"88050ca8",
   492 => x"0b80f4c4",
   493 => x"0b8c050c",
   494 => x"9f53a0a8",
   495 => x"5280f4d4",
   496 => x"518e933f",
   497 => x"9f53a0c8",
   498 => x"5280f6f0",
   499 => x"518e873f",
   500 => x"8a0bb2d8",
   501 => x"0ca3a851",
   502 => x"f9913fa0",
   503 => x"e851f98b",
   504 => x"3fa3a851",
   505 => x"f9853fa4",
   506 => x"d808802e",
   507 => x"83f138a1",
   508 => x"9851f8f7",
   509 => x"3fa3a851",
   510 => x"f8f13fa4",
   511 => x"d40852a1",
   512 => x"c451f8e7",
   513 => x"3fc808f8",
   514 => x"80110870",
   515 => x"a5f80c57",
   516 => x"55815880",
   517 => x"0ba4d408",
   518 => x"2582c538",
   519 => x"8c3d5b80",
   520 => x"c10b80f4",
   521 => x"f834810b",
   522 => x"80f7900c",
   523 => x"80c20b80",
   524 => x"f4fc3482",
   525 => x"5c835a9f",
   526 => x"53a1f452",
   527 => x"80f58051",
   528 => x"8d943f81",
   529 => x"5d800b80",
   530 => x"f5805380",
   531 => x"f6f05255",
   532 => x"86ed3f88",
   533 => x"08752e09",
   534 => x"81068338",
   535 => x"81557480",
   536 => x"f7900c7b",
   537 => x"70575574",
   538 => x"8325a038",
   539 => x"74101015",
   540 => x"fd055e8f",
   541 => x"3dfc0553",
   542 => x"83527551",
   543 => x"859d3f81",
   544 => x"1c705d70",
   545 => x"57558375",
   546 => x"24e2387d",
   547 => x"547453a5",
   548 => x"fc5280f5",
   549 => x"a8518593",
   550 => x"3f80f5a0",
   551 => x"08700857",
   552 => x"57b05376",
   553 => x"5275518c",
   554 => x"ad3f850b",
   555 => x"8c180c85",
   556 => x"0b8c170c",
   557 => x"7608760c",
   558 => x"80f5a008",
   559 => x"5574802e",
   560 => x"8a387408",
   561 => x"760c80f5",
   562 => x"a008558c",
   563 => x"155380f4",
   564 => x"f408528a",
   565 => x"5184c43f",
   566 => x"84160883",
   567 => x"a438860b",
   568 => x"8c170c88",
   569 => x"16528817",
   570 => x"085183cf",
   571 => x"3f80f5a0",
   572 => x"08700877",
   573 => x"0c558c16",
   574 => x"7054578a",
   575 => x"52760851",
   576 => x"84993f80",
   577 => x"c10b80f4",
   578 => x"fc335656",
   579 => x"757526a2",
   580 => x"3880c352",
   581 => x"755184fd",
   582 => x"3f88087d",
   583 => x"2e82b538",
   584 => x"81167081",
   585 => x"ff0680f4",
   586 => x"fc335757",
   587 => x"57747627",
   588 => x"e0387d7a",
   589 => x"7d293570",
   590 => x"5d8a1180",
   591 => x"f4f83380",
   592 => x"f4f4085a",
   593 => x"58515575",
   594 => x"80c12e82",
   595 => x"cc3878f7",
   596 => x"38811858",
   597 => x"a4d40878",
   598 => x"25fdc438",
   599 => x"a5f80856",
   600 => x"c808f880",
   601 => x"11087080",
   602 => x"f4bc0c70",
   603 => x"783170a5",
   604 => x"f40c54a2",
   605 => x"94535c5a",
   606 => x"f5f13fa5",
   607 => x"f4085680",
   608 => x"f7762580",
   609 => x"e038a4d4",
   610 => x"08707787",
   611 => x"e82935a5",
   612 => x"ec0c7671",
   613 => x"87e82935",
   614 => x"a5f00c76",
   615 => x"7184b929",
   616 => x"3580f5a4",
   617 => x"0c57a2a4",
   618 => x"51f5c03f",
   619 => x"a5ec0852",
   620 => x"a2d451f5",
   621 => x"b63fa2dc",
   622 => x"51f5b03f",
   623 => x"a5f00852",
   624 => x"a2d451f5",
   625 => x"a63f80f5",
   626 => x"a40852a3",
   627 => x"8c51f59b",
   628 => x"3fa3a851",
   629 => x"f5953f80",
   630 => x"0b880c8f",
   631 => x"3d0d04a3",
   632 => x"ac51fc8e",
   633 => x"39a3dc51",
   634 => x"f5813fa4",
   635 => x"9451f4fb",
   636 => x"3fa3a851",
   637 => x"f4f53fa5",
   638 => x"f408a4d4",
   639 => x"08707287",
   640 => x"e82935a5",
   641 => x"ec0c7171",
   642 => x"87e82935",
   643 => x"a5f00c71",
   644 => x"7184b929",
   645 => x"3580f5a4",
   646 => x"0c5856a2",
   647 => x"a451f4cb",
   648 => x"3fa5ec08",
   649 => x"52a2d451",
   650 => x"f4c13fa2",
   651 => x"dc51f4bb",
   652 => x"3fa5f008",
   653 => x"52a2d451",
   654 => x"f4b13f80",
   655 => x"f5a40852",
   656 => x"a38c51f4",
   657 => x"a63fa3a8",
   658 => x"51f4a03f",
   659 => x"800b880c",
   660 => x"8f3d0d04",
   661 => x"8f3df805",
   662 => x"52805180",
   663 => x"de3f9f53",
   664 => x"a4b45280",
   665 => x"f5805188",
   666 => x"ed3f7778",
   667 => x"80f4f40c",
   668 => x"81177081",
   669 => x"ff0680f4",
   670 => x"fc335858",
   671 => x"585afdad",
   672 => x"39760856",
   673 => x"b0537552",
   674 => x"765188ca",
   675 => x"3f80c10b",
   676 => x"80f4fc33",
   677 => x"5656fcf4",
   678 => x"39ff1570",
   679 => x"78317c0c",
   680 => x"598059fd",
   681 => x"ac39ff3d",
   682 => x"0d738232",
   683 => x"70307072",
   684 => x"07802588",
   685 => x"0c525283",
   686 => x"3d0d04fe",
   687 => x"3d0d7476",
   688 => x"71535452",
   689 => x"71822e83",
   690 => x"38835171",
   691 => x"812e9a38",
   692 => x"8172269f",
   693 => x"3871822e",
   694 => x"b8387184",
   695 => x"2ea93870",
   696 => x"730c7088",
   697 => x"0c843d0d",
   698 => x"0480e40b",
   699 => x"80f4f408",
   700 => x"258b3880",
   701 => x"730c7088",
   702 => x"0c843d0d",
   703 => x"0483730c",
   704 => x"70880c84",
   705 => x"3d0d0482",
   706 => x"730c7088",
   707 => x"0c843d0d",
   708 => x"0481730c",
   709 => x"70880c84",
   710 => x"3d0d0480",
   711 => x"3d0d7474",
   712 => x"14820571",
   713 => x"0c880c82",
   714 => x"3d0d04f7",
   715 => x"3d0d7b7d",
   716 => x"7f618512",
   717 => x"70822b75",
   718 => x"11707471",
   719 => x"70840553",
   720 => x"0c5a5a5d",
   721 => x"5b760c79",
   722 => x"80f8180c",
   723 => x"79861252",
   724 => x"57585a5a",
   725 => x"76762499",
   726 => x"3876b329",
   727 => x"822b7911",
   728 => x"51537673",
   729 => x"70840555",
   730 => x"0c811454",
   731 => x"757425f2",
   732 => x"387681cc",
   733 => x"2919fc11",
   734 => x"088105fc",
   735 => x"120c7a19",
   736 => x"70089fa0",
   737 => x"130c5856",
   738 => x"850b80f4",
   739 => x"f40c7588",
   740 => x"0c8b3d0d",
   741 => x"04fe3d0d",
   742 => x"02930533",
   743 => x"51800284",
   744 => x"05970533",
   745 => x"54527073",
   746 => x"2e883871",
   747 => x"880c843d",
   748 => x"0d047080",
   749 => x"f4f83481",
   750 => x"0b880c84",
   751 => x"3d0d04f8",
   752 => x"3d0d7a7c",
   753 => x"5956820b",
   754 => x"83195555",
   755 => x"74167033",
   756 => x"75335b51",
   757 => x"5372792e",
   758 => x"80c63880",
   759 => x"c10b8116",
   760 => x"81165656",
   761 => x"57827525",
   762 => x"e338ffa9",
   763 => x"177081ff",
   764 => x"06555973",
   765 => x"82268338",
   766 => x"87558153",
   767 => x"7680d22e",
   768 => x"98387752",
   769 => x"755186e7",
   770 => x"3f805372",
   771 => x"88082589",
   772 => x"38871580",
   773 => x"f4f40c81",
   774 => x"5372880c",
   775 => x"8a3d0d04",
   776 => x"7280f4f8",
   777 => x"34827525",
   778 => x"ffa238ff",
   779 => x"bd399408",
   780 => x"02940cfd",
   781 => x"3d0d8053",
   782 => x"94088c05",
   783 => x"08529408",
   784 => x"88050851",
   785 => x"82de3f88",
   786 => x"0870880c",
   787 => x"54853d0d",
   788 => x"940c0494",
   789 => x"0802940c",
   790 => x"fd3d0d81",
   791 => x"5394088c",
   792 => x"05085294",
   793 => x"08880508",
   794 => x"5182b93f",
   795 => x"88087088",
   796 => x"0c54853d",
   797 => x"0d940c04",
   798 => x"94080294",
   799 => x"0cf93d0d",
   800 => x"800b9408",
   801 => x"fc050c94",
   802 => x"08880508",
   803 => x"8025ab38",
   804 => x"94088805",
   805 => x"08309408",
   806 => x"88050c80",
   807 => x"0b9408f4",
   808 => x"050c9408",
   809 => x"fc050888",
   810 => x"38810b94",
   811 => x"08f4050c",
   812 => x"9408f405",
   813 => x"089408fc",
   814 => x"050c9408",
   815 => x"8c050880",
   816 => x"25ab3894",
   817 => x"088c0508",
   818 => x"3094088c",
   819 => x"050c800b",
   820 => x"9408f005",
   821 => x"0c9408fc",
   822 => x"05088838",
   823 => x"810b9408",
   824 => x"f0050c94",
   825 => x"08f00508",
   826 => x"9408fc05",
   827 => x"0c805394",
   828 => x"088c0508",
   829 => x"52940888",
   830 => x"05085181",
   831 => x"a73f8808",
   832 => x"709408f8",
   833 => x"050c5494",
   834 => x"08fc0508",
   835 => x"802e8c38",
   836 => x"9408f805",
   837 => x"08309408",
   838 => x"f8050c94",
   839 => x"08f80508",
   840 => x"70880c54",
   841 => x"893d0d94",
   842 => x"0c049408",
   843 => x"02940cfb",
   844 => x"3d0d800b",
   845 => x"9408fc05",
   846 => x"0c940888",
   847 => x"05088025",
   848 => x"93389408",
   849 => x"88050830",
   850 => x"94088805",
   851 => x"0c810b94",
   852 => x"08fc050c",
   853 => x"94088c05",
   854 => x"0880258c",
   855 => x"3894088c",
   856 => x"05083094",
   857 => x"088c050c",
   858 => x"81539408",
   859 => x"8c050852",
   860 => x"94088805",
   861 => x"0851ad3f",
   862 => x"88087094",
   863 => x"08f8050c",
   864 => x"549408fc",
   865 => x"0508802e",
   866 => x"8c389408",
   867 => x"f8050830",
   868 => x"9408f805",
   869 => x"0c9408f8",
   870 => x"05087088",
   871 => x"0c54873d",
   872 => x"0d940c04",
   873 => x"94080294",
   874 => x"0cfd3d0d",
   875 => x"810b9408",
   876 => x"fc050c80",
   877 => x"0b9408f8",
   878 => x"050c9408",
   879 => x"8c050894",
   880 => x"08880508",
   881 => x"27ac3894",
   882 => x"08fc0508",
   883 => x"802ea338",
   884 => x"800b9408",
   885 => x"8c050824",
   886 => x"99389408",
   887 => x"8c050810",
   888 => x"94088c05",
   889 => x"0c9408fc",
   890 => x"05081094",
   891 => x"08fc050c",
   892 => x"c9399408",
   893 => x"fc050880",
   894 => x"2e80c938",
   895 => x"94088c05",
   896 => x"08940888",
   897 => x"050826a1",
   898 => x"38940888",
   899 => x"05089408",
   900 => x"8c050831",
   901 => x"94088805",
   902 => x"0c9408f8",
   903 => x"05089408",
   904 => x"fc050807",
   905 => x"9408f805",
   906 => x"0c9408fc",
   907 => x"0508812a",
   908 => x"9408fc05",
   909 => x"0c94088c",
   910 => x"0508812a",
   911 => x"94088c05",
   912 => x"0cffaf39",
   913 => x"94089005",
   914 => x"08802e8f",
   915 => x"38940888",
   916 => x"05087094",
   917 => x"08f4050c",
   918 => x"518d3994",
   919 => x"08f80508",
   920 => x"709408f4",
   921 => x"050c5194",
   922 => x"08f40508",
   923 => x"880c853d",
   924 => x"0d940c04",
   925 => x"94080294",
   926 => x"0cff3d0d",
   927 => x"800b9408",
   928 => x"fc050c94",
   929 => x"08880508",
   930 => x"8106ff11",
   931 => x"70097094",
   932 => x"088c0508",
   933 => x"069408fc",
   934 => x"05081194",
   935 => x"08fc050c",
   936 => x"94088805",
   937 => x"08812a94",
   938 => x"0888050c",
   939 => x"94088c05",
   940 => x"08109408",
   941 => x"8c050c51",
   942 => x"51515194",
   943 => x"08880508",
   944 => x"802e8438",
   945 => x"ffbd3994",
   946 => x"08fc0508",
   947 => x"70880c51",
   948 => x"833d0d94",
   949 => x"0c04fc3d",
   950 => x"0d767079",
   951 => x"7b555555",
   952 => x"558f7227",
   953 => x"8c387275",
   954 => x"07830651",
   955 => x"70802ea7",
   956 => x"38ff1252",
   957 => x"71ff2e98",
   958 => x"38727081",
   959 => x"05543374",
   960 => x"70810556",
   961 => x"34ff1252",
   962 => x"71ff2e09",
   963 => x"8106ea38",
   964 => x"74880c86",
   965 => x"3d0d0474",
   966 => x"51727084",
   967 => x"05540871",
   968 => x"70840553",
   969 => x"0c727084",
   970 => x"05540871",
   971 => x"70840553",
   972 => x"0c727084",
   973 => x"05540871",
   974 => x"70840553",
   975 => x"0c727084",
   976 => x"05540871",
   977 => x"70840553",
   978 => x"0cf01252",
   979 => x"718f26c9",
   980 => x"38837227",
   981 => x"95387270",
   982 => x"84055408",
   983 => x"71708405",
   984 => x"530cfc12",
   985 => x"52718326",
   986 => x"ed387054",
   987 => x"ff8339fb",
   988 => x"3d0d7779",
   989 => x"70720783",
   990 => x"06535452",
   991 => x"70933871",
   992 => x"73730854",
   993 => x"56547173",
   994 => x"082e80c4",
   995 => x"38737554",
   996 => x"52713370",
   997 => x"81ff0652",
   998 => x"5470802e",
   999 => x"9d387233",
  1000 => x"5570752e",
  1001 => x"09810695",
  1002 => x"38811281",
  1003 => x"14713370",
  1004 => x"81ff0654",
  1005 => x"56545270",
  1006 => x"e5387233",
  1007 => x"557381ff",
  1008 => x"067581ff",
  1009 => x"06717131",
  1010 => x"880c5252",
  1011 => x"873d0d04",
  1012 => x"710970f7",
  1013 => x"fbfdff14",
  1014 => x"0670f884",
  1015 => x"82818006",
  1016 => x"51515170",
  1017 => x"97388414",
  1018 => x"84167108",
  1019 => x"54565471",
  1020 => x"75082edc",
  1021 => x"38737554",
  1022 => x"52ff9639",
  1023 => x"800b880c",
  1024 => x"873d0d04",
  1025 => x"00ffffff",
  1026 => x"ff00ffff",
  1027 => x"ffff00ff",
  1028 => x"ffffff00",
  1029 => x"30313233",
  1030 => x"34353637",
  1031 => x"38394142",
  1032 => x"43444546",
  1033 => x"00000000",
  1034 => x"44485259",
  1035 => x"53544f4e",
  1036 => x"45205052",
  1037 => x"4f475241",
  1038 => x"4d2c2053",
  1039 => x"4f4d4520",
  1040 => x"53545249",
  1041 => x"4e470000",
  1042 => x"44485259",
  1043 => x"53544f4e",
  1044 => x"45205052",
  1045 => x"4f475241",
  1046 => x"4d2c2031",
  1047 => x"27535420",
  1048 => x"53545249",
  1049 => x"4e470000",
  1050 => x"44687279",
  1051 => x"73746f6e",
  1052 => x"65204265",
  1053 => x"6e63686d",
  1054 => x"61726b2c",
  1055 => x"20566572",
  1056 => x"73696f6e",
  1057 => x"20322e31",
  1058 => x"20284c61",
  1059 => x"6e677561",
  1060 => x"67653a20",
  1061 => x"43290a00",
  1062 => x"50726f67",
  1063 => x"72616d20",
  1064 => x"636f6d70",
  1065 => x"696c6564",
  1066 => x"20776974",
  1067 => x"68202772",
  1068 => x"65676973",
  1069 => x"74657227",
  1070 => x"20617474",
  1071 => x"72696275",
  1072 => x"74650a00",
  1073 => x"45786563",
  1074 => x"7574696f",
  1075 => x"6e207374",
  1076 => x"61727473",
  1077 => x"2c202564",
  1078 => x"2072756e",
  1079 => x"73207468",
  1080 => x"726f7567",
  1081 => x"68204468",
  1082 => x"72797374",
  1083 => x"6f6e650a",
  1084 => x"00000000",
  1085 => x"44485259",
  1086 => x"53544f4e",
  1087 => x"45205052",
  1088 => x"4f475241",
  1089 => x"4d2c2032",
  1090 => x"274e4420",
  1091 => x"53545249",
  1092 => x"4e470000",
  1093 => x"55736572",
  1094 => x"2074696d",
  1095 => x"653a2025",
  1096 => x"640a0000",
  1097 => x"4d696372",
  1098 => x"6f736563",
  1099 => x"6f6e6473",
  1100 => x"20666f72",
  1101 => x"206f6e65",
  1102 => x"2072756e",
  1103 => x"20746872",
  1104 => x"6f756768",
  1105 => x"20446872",
  1106 => x"7973746f",
  1107 => x"6e653a20",
  1108 => x"00000000",
  1109 => x"2564200a",
  1110 => x"00000000",
  1111 => x"44687279",
  1112 => x"73746f6e",
  1113 => x"65732070",
  1114 => x"65722053",
  1115 => x"65636f6e",
  1116 => x"643a2020",
  1117 => x"20202020",
  1118 => x"20202020",
  1119 => x"20202020",
  1120 => x"20202020",
  1121 => x"20202020",
  1122 => x"00000000",
  1123 => x"56415820",
  1124 => x"4d495053",
  1125 => x"20726174",
  1126 => x"696e6720",
  1127 => x"2a203130",
  1128 => x"3030203d",
  1129 => x"20256420",
  1130 => x"0a000000",
  1131 => x"50726f67",
  1132 => x"72616d20",
  1133 => x"636f6d70",
  1134 => x"696c6564",
  1135 => x"20776974",
  1136 => x"686f7574",
  1137 => x"20277265",
  1138 => x"67697374",
  1139 => x"65722720",
  1140 => x"61747472",
  1141 => x"69627574",
  1142 => x"650a0000",
  1143 => x"4d656173",
  1144 => x"75726564",
  1145 => x"2074696d",
  1146 => x"6520746f",
  1147 => x"6f20736d",
  1148 => x"616c6c20",
  1149 => x"746f206f",
  1150 => x"62746169",
  1151 => x"6e206d65",
  1152 => x"616e696e",
  1153 => x"6766756c",
  1154 => x"20726573",
  1155 => x"756c7473",
  1156 => x"0a000000",
  1157 => x"506c6561",
  1158 => x"73652069",
  1159 => x"6e637265",
  1160 => x"61736520",
  1161 => x"6e756d62",
  1162 => x"6572206f",
  1163 => x"66207275",
  1164 => x"6e730a00",
  1165 => x"44485259",
  1166 => x"53544f4e",
  1167 => x"45205052",
  1168 => x"4f475241",
  1169 => x"4d2c2033",
  1170 => x"27524420",
  1171 => x"53545249",
  1172 => x"4e470000",
  1173 => x"000061a8",
  1174 => x"00000000",
	others => x"00000000"
);

begin

process (clk)
begin
	if (clk'event and clk = '1') then
		if (from_zpu.memAWriteEnable = '1') and (from_zpu.memBWriteEnable = '1') and (from_zpu.memAAddr=from_zpu.memBAddr) and (from_zpu.memAWrite/=from_zpu.memBWrite) then
			report "write collision" severity failure;
		end if;
	
		if (from_zpu.memAWriteEnable = '1') then
			ram(to_integer(unsigned(from_zpu.memAAddr(maxAddrBitBRAM downto 2)))) := from_zpu.memAWrite;
			to_zpu.memARead <= from_zpu.memAWrite;
		else
			to_zpu.memARead <= ram(to_integer(unsigned(from_zpu.memAAddr(maxAddrBitBRAM downto 2))));
		end if;
	end if;
end process;

process (clk)
begin
	if (clk'event and clk = '1') then
		if (from_zpu.memBWriteEnable = '1') then
			ram(to_integer(unsigned(from_zpu.memBAddr(maxAddrBitBRAM downto 2)))) := from_zpu.memBWrite;
			to_zpu.memBRead <= from_zpu.memBWrite;
		else
			to_zpu.memBRead <= ram(to_integer(unsigned(from_zpu.memBAddr(maxAddrBitBRAM downto 2))));
		end if;
	end if;
end process;


end arch;

