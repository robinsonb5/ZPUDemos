-- ZPU
--
-- Copyright 2004-2008 oharboe - �yvind Harboe - oyvind.harboe@zylin.com
-- Modified by Alastair M. Robinson for the ZPUFlex project.
--
-- The FreeBSD license
-- 
-- Redistribution and use in source and binary forms, with or without
-- modification, are permitted provided that the following conditions
-- are met:
-- 
-- 1. Redistributions of source code must retain the above copyright
--    notice, this list of conditions and the following disclaimer.
-- 2. Redistributions in binary form must reproduce the above
--    copyright notice, this list of conditions and the following
--    disclaimer in the documentation and/or other materials
--    provided with the distribution.
-- 
-- THIS SOFTWARE IS PROVIDED BY THE ZPU PROJECT ``AS IS'' AND ANY
-- EXPRESS OR IMPLIED WARRANTIES, INCLUDING, BUT NOT LIMITED TO,
-- THE IMPLIED WARRANTIES OF MERCHANTABILITY AND FITNESS FOR A
-- PARTICULAR PURPOSE ARE DISCLAIMED. IN NO EVENT SHALL THE
-- ZPU PROJECT OR CONTRIBUTORS BE LIABLE FOR ANY DIRECT,
-- INDIRECT, INCIDENTAL, SPECIAL, EXEMPLARY, OR CONSEQUENTIAL DAMAGES
-- (INCLUDING, BUT NOT LIMITED TO, PROCUREMENT OF SUBSTITUTE GOODS
-- OR SERVICES; LOSS OF USE, DATA, OR PROFITS; OR BUSINESS INTERRUPTION)
-- HOWEVER CAUSED AND ON ANY THEORY OF LIABILITY, WHETHER IN CONTRACT,
-- STRICT LIABILITY, OR TORT (INCLUDING NEGLIGENCE OR OTHERWISE)
-- ARISING IN ANY WAY OUT OF THE USE OF THIS SOFTWARE, EVEN IF
-- ADVISED OF THE POSSIBILITY OF SUCH DAMAGE.
-- 
-- The views and conclusions contained in the software and documentation
-- are those of the authors and should not be interpreted as representing
-- official policies, either expressed or implied, of the ZPU Project.

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;


library work;
use work.zpu_config.all;
use work.zpupkg.all;

entity SDRAMTest_ROM is
generic
	(
		maxAddrBitBRAM : integer := maxAddrBitBRAMLimit -- Specify your actual ROM size to save LEs and unnecessary block RAM usage.
	);
port (
	clk : in std_logic;
	areset : in std_logic := '0';
	from_zpu : in ZPU_ToROM;
	to_zpu : out ZPU_FromROM
);
end SDRAMTest_ROM;

architecture arch of SDRAMTest_ROM is

type ram_type is array(natural range 0 to ((2**(maxAddrBitBRAM+1))/4)-1) of std_logic_vector(wordSize-1 downto 0);

shared variable ram : ram_type :=
(
     0 => x"84808080",
     1 => x"ed040000",
     2 => x"00000000",
     3 => x"84808080",
     4 => x"880d8004",
     5 => x"84808080",
     6 => x"940471fd",
     7 => x"06087283",
     8 => x"06098105",
     9 => x"8205832b",
    10 => x"2a83ffff",
    11 => x"06520471",
    12 => x"fc060872",
    13 => x"83060981",
    14 => x"05830510",
    15 => x"10102a81",
    16 => x"ff065204",
    17 => x"71fc0608",
    18 => x"8480808f",
    19 => x"dc738306",
    20 => x"10100508",
    21 => x"067381ff",
    22 => x"06738306",
    23 => x"09810583",
    24 => x"05101010",
    25 => x"2b0772fc",
    26 => x"060c5151",
    27 => x"04028405",
    28 => x"84808080",
    29 => x"880c8480",
    30 => x"8080940b",
    31 => x"8480808c",
    32 => x"c9040000",
    33 => x"02c0050d",
    34 => x"0280c405",
    35 => x"84808096",
    36 => x"c85c5c80",
    37 => x"7c708405",
    38 => x"5e08715f",
    39 => x"5f587d70",
    40 => x"84055f08",
    41 => x"57805a76",
    42 => x"982a7788",
    43 => x"2b585574",
    44 => x"802e82a3",
    45 => x"387c802e",
    46 => x"80c53880",
    47 => x"5d7480e4",
    48 => x"2e81bb38",
    49 => x"7480e426",
    50 => x"80f13874",
    51 => x"80e32e80",
    52 => x"c838a551",
    53 => x"84808083",
    54 => x"f92d7451",
    55 => x"84808083",
    56 => x"f92d8218",
    57 => x"58811a5a",
    58 => x"837a25ff",
    59 => x"ba3874ff",
    60 => x"ad387e84",
    61 => x"808095e8",
    62 => x"0c0280c0",
    63 => x"050d0474",
    64 => x"a52e0981",
    65 => x"069b3881",
    66 => x"0b811b5b",
    67 => x"5d837a25",
    68 => x"ff953884",
    69 => x"808081ee",
    70 => x"047b841d",
    71 => x"7108575d",
    72 => x"54745184",
    73 => x"808083f9",
    74 => x"2d811881",
    75 => x"1b5b5883",
    76 => x"7a25fef3",
    77 => x"38848080",
    78 => x"81ee0474",
    79 => x"80f32e09",
    80 => x"8106ff8e",
    81 => x"387b841d",
    82 => x"71087054",
    83 => x"5d5d5384",
    84 => x"8080849e",
    85 => x"2d800bff",
    86 => x"11545280",
    87 => x"7225ff85",
    88 => x"387a7081",
    89 => x"055c3370",
    90 => x"52558480",
    91 => x"8083f92d",
    92 => x"811873ff",
    93 => x"15555358",
    94 => x"84808082",
    95 => x"db047b84",
    96 => x"1d71087f",
    97 => x"5c565d52",
    98 => x"80742480",
    99 => x"d7388756",
   100 => x"739c2a74",
   101 => x"842b5552",
   102 => x"71802e83",
   103 => x"388159b7",
   104 => x"12537189",
   105 => x"248438b0",
   106 => x"12537895",
   107 => x"38ff1656",
   108 => x"758025dc",
   109 => x"38800bff",
   110 => x"11545284",
   111 => x"808082db",
   112 => x"04725184",
   113 => x"808083f9",
   114 => x"2dff1656",
   115 => x"758025c0",
   116 => x"38848080",
   117 => x"83b50477",
   118 => x"84808095",
   119 => x"e80c0280",
   120 => x"c0050d04",
   121 => x"ad518480",
   122 => x"8083f92d",
   123 => x"73098105",
   124 => x"54875684",
   125 => x"80808390",
   126 => x"0402f805",
   127 => x"0d7352c0",
   128 => x"0870882a",
   129 => x"70810651",
   130 => x"51517080",
   131 => x"2ef13871",
   132 => x"c00c7184",
   133 => x"808095e8",
   134 => x"0c028805",
   135 => x"0d0402e8",
   136 => x"050d8078",
   137 => x"57557570",
   138 => x"84055708",
   139 => x"53805472",
   140 => x"982a7388",
   141 => x"2b545271",
   142 => x"802ea238",
   143 => x"c0087088",
   144 => x"2a708106",
   145 => x"51515170",
   146 => x"802ef138",
   147 => x"71c00c81",
   148 => x"15811555",
   149 => x"55837425",
   150 => x"d63871ca",
   151 => x"38748480",
   152 => x"8095e80c",
   153 => x"0298050d",
   154 => x"0402f405",
   155 => x"0d747652",
   156 => x"53807125",
   157 => x"90387052",
   158 => x"72708405",
   159 => x"5408ff13",
   160 => x"535171f4",
   161 => x"38028c05",
   162 => x"0d0402d4",
   163 => x"050d7c7e",
   164 => x"5c58810b",
   165 => x"8480808f",
   166 => x"ec585a83",
   167 => x"59760878",
   168 => x"0c770877",
   169 => x"08565473",
   170 => x"752e9438",
   171 => x"77085374",
   172 => x"52848080",
   173 => x"8ffc5184",
   174 => x"80808184",
   175 => x"2d805a77",
   176 => x"56807b25",
   177 => x"90387a55",
   178 => x"75708405",
   179 => x"5708ff16",
   180 => x"565474f4",
   181 => x"38770877",
   182 => x"08565675",
   183 => x"752e9438",
   184 => x"77085374",
   185 => x"52848080",
   186 => x"90bc5184",
   187 => x"80808184",
   188 => x"2d805aff",
   189 => x"19841858",
   190 => x"59788025",
   191 => x"ff9f3879",
   192 => x"84808095",
   193 => x"e80c02ac",
   194 => x"050d0402",
   195 => x"e4050d78",
   196 => x"7a555681",
   197 => x"5785aad5",
   198 => x"aad5760c",
   199 => x"fad5aad5",
   200 => x"aa0b8c17",
   201 => x"0ccc7634",
   202 => x"b30b8f17",
   203 => x"34750853",
   204 => x"72fce2d5",
   205 => x"aad52e92",
   206 => x"38750852",
   207 => x"84808090",
   208 => x"fc518480",
   209 => x"8081842d",
   210 => x"80578c16",
   211 => x"085574fa",
   212 => x"d5aad4b3",
   213 => x"2e93388c",
   214 => x"16085284",
   215 => x"808091b8",
   216 => x"51848080",
   217 => x"81842d80",
   218 => x"57755580",
   219 => x"74258e38",
   220 => x"74708405",
   221 => x"5608ff15",
   222 => x"555373f4",
   223 => x"38750854",
   224 => x"73fce2d5",
   225 => x"aad52e92",
   226 => x"38750852",
   227 => x"84808091",
   228 => x"f4518480",
   229 => x"8081842d",
   230 => x"80578c16",
   231 => x"085372fa",
   232 => x"d5aad4b3",
   233 => x"2e93388c",
   234 => x"16085284",
   235 => x"808092b0",
   236 => x"51848080",
   237 => x"81842d80",
   238 => x"57768480",
   239 => x"8095e80c",
   240 => x"029c050d",
   241 => x"0402c405",
   242 => x"0d605b80",
   243 => x"62908080",
   244 => x"29ff0584",
   245 => x"808092ec",
   246 => x"53405a84",
   247 => x"80808184",
   248 => x"2d80e1b3",
   249 => x"5780fe5e",
   250 => x"ae518480",
   251 => x"8083f92d",
   252 => x"76107096",
   253 => x"2a810656",
   254 => x"5774802e",
   255 => x"85387681",
   256 => x"07577695",
   257 => x"2a810658",
   258 => x"77802e85",
   259 => x"38768132",
   260 => x"57787707",
   261 => x"7f06775e",
   262 => x"598fffff",
   263 => x"5876bfff",
   264 => x"ff06707a",
   265 => x"32822b7c",
   266 => x"11515776",
   267 => x"0c761070",
   268 => x"962a8106",
   269 => x"56577480",
   270 => x"2e853876",
   271 => x"81075776",
   272 => x"952a8106",
   273 => x"5574802e",
   274 => x"85387681",
   275 => x"3257ff18",
   276 => x"58778025",
   277 => x"c8387c57",
   278 => x"8fffff58",
   279 => x"76bfffff",
   280 => x"06707a32",
   281 => x"822b7c05",
   282 => x"7008575e",
   283 => x"5674762e",
   284 => x"80ea3880",
   285 => x"7a538480",
   286 => x"8092fc52",
   287 => x"5c848080",
   288 => x"81842d74",
   289 => x"54755375",
   290 => x"52848080",
   291 => x"93905184",
   292 => x"80808184",
   293 => x"2d7b5a76",
   294 => x"1070962a",
   295 => x"81065757",
   296 => x"75802e85",
   297 => x"38768107",
   298 => x"5776952a",
   299 => x"81065574",
   300 => x"802e8538",
   301 => x"76813257",
   302 => x"ff185877",
   303 => x"8025ff9c",
   304 => x"38ff1e5e",
   305 => x"7dfea138",
   306 => x"8a518480",
   307 => x"8083f92d",
   308 => x"7b848080",
   309 => x"95e80c02",
   310 => x"bc050d04",
   311 => x"811a5a84",
   312 => x"80808997",
   313 => x"0402cc05",
   314 => x"0d7e605e",
   315 => x"58815a80",
   316 => x"5b80c07a",
   317 => x"585c85ad",
   318 => x"a989bb78",
   319 => x"0c795981",
   320 => x"56975576",
   321 => x"7607822b",
   322 => x"78115154",
   323 => x"85ada989",
   324 => x"bb740c75",
   325 => x"10ff1656",
   326 => x"56748025",
   327 => x"e6387610",
   328 => x"811a5a57",
   329 => x"987925d7",
   330 => x"38775680",
   331 => x"7d259038",
   332 => x"7c557570",
   333 => x"84055708",
   334 => x"ff165654",
   335 => x"74f43881",
   336 => x"57ff8787",
   337 => x"a5c3780c",
   338 => x"97597682",
   339 => x"2b781170",
   340 => x"085f5656",
   341 => x"7cff8787",
   342 => x"a5c32e80",
   343 => x"cc387408",
   344 => x"547385ad",
   345 => x"a989bb2e",
   346 => x"94388075",
   347 => x"08547653",
   348 => x"84808093",
   349 => x"b8525a84",
   350 => x"80808184",
   351 => x"2d7610ff",
   352 => x"1a5a5778",
   353 => x"8025c338",
   354 => x"7a822b56",
   355 => x"75b1387b",
   356 => x"52848080",
   357 => x"93d85184",
   358 => x"80808184",
   359 => x"2d7b8480",
   360 => x"8095e80c",
   361 => x"02b4050d",
   362 => x"047a7707",
   363 => x"7710ff1b",
   364 => x"5b585b78",
   365 => x"8025ff92",
   366 => x"38848080",
   367 => x"8b880475",
   368 => x"52848080",
   369 => x"94945184",
   370 => x"80808184",
   371 => x"2d75992a",
   372 => x"81328106",
   373 => x"70098105",
   374 => x"71077009",
   375 => x"709f2c7d",
   376 => x"0679109f",
   377 => x"fffffc06",
   378 => x"60812a41",
   379 => x"5a5d5758",
   380 => x"5975da38",
   381 => x"79098105",
   382 => x"707b079f",
   383 => x"2a55567b",
   384 => x"bf268438",
   385 => x"739d3881",
   386 => x"70538480",
   387 => x"8093d852",
   388 => x"5c848080",
   389 => x"81842d7b",
   390 => x"84808095",
   391 => x"e80c02b4",
   392 => x"050d0484",
   393 => x"808094ac",
   394 => x"51848080",
   395 => x"81842d7b",
   396 => x"52848080",
   397 => x"93d85184",
   398 => x"80808184",
   399 => x"2d7b8480",
   400 => x"8095e80c",
   401 => x"02b4050d",
   402 => x"0402dc05",
   403 => x"0d810b84",
   404 => x"80808fec",
   405 => x"58588359",
   406 => x"7608800c",
   407 => x"80087708",
   408 => x"56547375",
   409 => x"2e943880",
   410 => x"08537452",
   411 => x"8480808f",
   412 => x"fc518480",
   413 => x"8081842d",
   414 => x"80588070",
   415 => x"57557570",
   416 => x"84055708",
   417 => x"81165654",
   418 => x"a0807524",
   419 => x"f1388008",
   420 => x"77085656",
   421 => x"75752e94",
   422 => x"38800853",
   423 => x"74528480",
   424 => x"8090bc51",
   425 => x"84808081",
   426 => x"842d8058",
   427 => x"ff198418",
   428 => x"58597880",
   429 => x"25ffa138",
   430 => x"77802e8d",
   431 => x"38848080",
   432 => x"94f85184",
   433 => x"80808184",
   434 => x"2d815785",
   435 => x"aad5aad5",
   436 => x"0b800cfa",
   437 => x"d5aad5aa",
   438 => x"0b8c0ccc",
   439 => x"0b8034b3",
   440 => x"0b8f3480",
   441 => x"085574fc",
   442 => x"e2d5aad5",
   443 => x"2e923880",
   444 => x"08528480",
   445 => x"8090fc51",
   446 => x"84808081",
   447 => x"842d8057",
   448 => x"8c085877",
   449 => x"fad5aad4",
   450 => x"b32e9238",
   451 => x"8c085284",
   452 => x"808091b8",
   453 => x"51848080",
   454 => x"81842d80",
   455 => x"57807057",
   456 => x"55757084",
   457 => x"05570881",
   458 => x"165654a0",
   459 => x"807524f1",
   460 => x"38800859",
   461 => x"78fce2d5",
   462 => x"aad52e92",
   463 => x"38800852",
   464 => x"84808091",
   465 => x"f4518480",
   466 => x"8081842d",
   467 => x"80578c08",
   468 => x"5473fad5",
   469 => x"aad4b32e",
   470 => x"80ea388c",
   471 => x"08528480",
   472 => x"8092b051",
   473 => x"84808081",
   474 => x"842da080",
   475 => x"52805184",
   476 => x"808089e5",
   477 => x"2d848080",
   478 => x"95e80854",
   479 => x"84808095",
   480 => x"e808802e",
   481 => x"8d388480",
   482 => x"80959c51",
   483 => x"84808081",
   484 => x"842d7352",
   485 => x"80518480",
   486 => x"8087c52d",
   487 => x"84808095",
   488 => x"e808802e",
   489 => x"fda73884",
   490 => x"808095b4",
   491 => x"51848080",
   492 => x"81842d81",
   493 => x"0b848080",
   494 => x"8fec5858",
   495 => x"83598480",
   496 => x"808cd804",
   497 => x"76802eff",
   498 => x"a1388480",
   499 => x"8095cc51",
   500 => x"84808081",
   501 => x"842d8480",
   502 => x"808eea04",
   503 => x"00ffffff",
   504 => x"ff00ffff",
   505 => x"ffff00ff",
   506 => x"ffffff00",
   507 => x"00000000",
   508 => x"55555555",
   509 => x"aaaaaaaa",
   510 => x"ffffffff",
   511 => x"53616e69",
   512 => x"74792063",
   513 => x"6865636b",
   514 => x"20666169",
   515 => x"6c656420",
   516 => x"28626566",
   517 => x"6f726520",
   518 => x"63616368",
   519 => x"65207265",
   520 => x"66726573",
   521 => x"6829206f",
   522 => x"6e203078",
   523 => x"25642028",
   524 => x"676f7420",
   525 => x"30782564",
   526 => x"290a0000",
   527 => x"53616e69",
   528 => x"74792063",
   529 => x"6865636b",
   530 => x"20666169",
   531 => x"6c656420",
   532 => x"28616674",
   533 => x"65722063",
   534 => x"61636865",
   535 => x"20726566",
   536 => x"72657368",
   537 => x"29206f6e",
   538 => x"20307825",
   539 => x"64202867",
   540 => x"6f742030",
   541 => x"78256429",
   542 => x"0a000000",
   543 => x"42797465",
   544 => x"20636865",
   545 => x"636b2066",
   546 => x"61696c65",
   547 => x"64202862",
   548 => x"65666f72",
   549 => x"65206361",
   550 => x"63686520",
   551 => x"72656672",
   552 => x"65736829",
   553 => x"20617420",
   554 => x"30202867",
   555 => x"6f742030",
   556 => x"78256429",
   557 => x"0a000000",
   558 => x"42797465",
   559 => x"20636865",
   560 => x"636b2066",
   561 => x"61696c65",
   562 => x"64202862",
   563 => x"65666f72",
   564 => x"65206361",
   565 => x"63686520",
   566 => x"72656672",
   567 => x"65736829",
   568 => x"20617420",
   569 => x"33202867",
   570 => x"6f742030",
   571 => x"78256429",
   572 => x"0a000000",
   573 => x"42797465",
   574 => x"20636865",
   575 => x"636b2066",
   576 => x"61696c65",
   577 => x"64202861",
   578 => x"66746572",
   579 => x"20636163",
   580 => x"68652072",
   581 => x"65667265",
   582 => x"73682920",
   583 => x"61742030",
   584 => x"2028676f",
   585 => x"74203078",
   586 => x"2564290a",
   587 => x"00000000",
   588 => x"42797465",
   589 => x"20636865",
   590 => x"636b2066",
   591 => x"61696c65",
   592 => x"64202861",
   593 => x"66746572",
   594 => x"20636163",
   595 => x"68652072",
   596 => x"65667265",
   597 => x"73682920",
   598 => x"61742033",
   599 => x"2028676f",
   600 => x"74203078",
   601 => x"2564290a",
   602 => x"00000000",
   603 => x"43686563",
   604 => x"6b696e67",
   605 => x"206d656d",
   606 => x"6f727900",
   607 => x"30782564",
   608 => x"20676f6f",
   609 => x"64207265",
   610 => x"6164732c",
   611 => x"20000000",
   612 => x"4572726f",
   613 => x"72206174",
   614 => x"20307825",
   615 => x"642c2065",
   616 => x"78706563",
   617 => x"74656420",
   618 => x"30782564",
   619 => x"2c20676f",
   620 => x"74203078",
   621 => x"25640a00",
   622 => x"42616420",
   623 => x"64617461",
   624 => x"20666f75",
   625 => x"6e642061",
   626 => x"74203078",
   627 => x"25642028",
   628 => x"30782564",
   629 => x"290a0000",
   630 => x"53445241",
   631 => x"4d207369",
   632 => x"7a652028",
   633 => x"61737375",
   634 => x"6d696e67",
   635 => x"206e6f20",
   636 => x"61646472",
   637 => x"65737320",
   638 => x"6661756c",
   639 => x"74732920",
   640 => x"69732030",
   641 => x"78256420",
   642 => x"6d656761",
   643 => x"62797465",
   644 => x"730a0000",
   645 => x"416c6961",
   646 => x"73657320",
   647 => x"666f756e",
   648 => x"64206174",
   649 => x"20307825",
   650 => x"640a0000",
   651 => x"28416c69",
   652 => x"61736573",
   653 => x"2070726f",
   654 => x"6261626c",
   655 => x"79207369",
   656 => x"6d706c79",
   657 => x"20696e64",
   658 => x"69636174",
   659 => x"65207468",
   660 => x"61742052",
   661 => x"414d0a69",
   662 => x"7320736d",
   663 => x"616c6c65",
   664 => x"72207468",
   665 => x"616e2036",
   666 => x"34206d65",
   667 => x"67616279",
   668 => x"74657329",
   669 => x"0a000000",
   670 => x"46697273",
   671 => x"74207374",
   672 => x"61676520",
   673 => x"73616e69",
   674 => x"74792063",
   675 => x"6865636b",
   676 => x"20706173",
   677 => x"7365642e",
   678 => x"0a000000",
   679 => x"41646472",
   680 => x"65737320",
   681 => x"63686563",
   682 => x"6b207061",
   683 => x"73736564",
   684 => x"2e0a0000",
   685 => x"4c465352",
   686 => x"20636865",
   687 => x"636b2070",
   688 => x"61737365",
   689 => x"642e0a0a",
   690 => x"00000000",
   691 => x"42797465",
   692 => x"20286471",
   693 => x"6d292063",
   694 => x"6865636b",
   695 => x"20706173",
   696 => x"7365640a",
   697 => x"00000000",
	others => x"00000000"
);

begin

process (clk)
begin
	if (clk'event and clk = '1') then
		if (from_zpu.memAWriteEnable = '1') and (from_zpu.memBWriteEnable = '1') and (from_zpu.memAAddr=from_zpu.memBAddr) and (from_zpu.memAWrite/=from_zpu.memBWrite) then
			report "write collision" severity failure;
		end if;
	
		if (from_zpu.memAWriteEnable = '1') then
			ram(to_integer(unsigned(from_zpu.memAAddr(maxAddrBitBRAM downto 2)))) := from_zpu.memAWrite;
			to_zpu.memARead <= from_zpu.memAWrite;
		else
			to_zpu.memARead <= ram(to_integer(unsigned(from_zpu.memAAddr(maxAddrBitBRAM downto 2))));
		end if;
	end if;
end process;

process (clk)
begin
	if (clk'event and clk = '1') then
		if (from_zpu.memBWriteEnable = '1') then
			ram(to_integer(unsigned(from_zpu.memBAddr(maxAddrBitBRAM downto 2)))) := from_zpu.memBWrite;
			to_zpu.memBRead <= from_zpu.memBWrite;
		else
			to_zpu.memBRead <= ram(to_integer(unsigned(from_zpu.memBAddr(maxAddrBitBRAM downto 2))));
		end if;
	end if;
end process;


end arch;

