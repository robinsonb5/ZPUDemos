-- ZPU
--
-- Copyright 2004-2008 oharboe - �yvind Harboe - oyvind.harboe@zylin.com
-- Modified by Alastair M. Robinson for the ZPUFlex project.
--
-- The FreeBSD license
-- 
-- Redistribution and use in source and binary forms, with or without
-- modification, are permitted provided that the following conditions
-- are met:
-- 
-- 1. Redistributions of source code must retain the above copyright
--    notice, this list of conditions and the following disclaimer.
-- 2. Redistributions in binary form must reproduce the above
--    copyright notice, this list of conditions and the following
--    disclaimer in the documentation and/or other materials
--    provided with the distribution.
-- 
-- THIS SOFTWARE IS PROVIDED BY THE ZPU PROJECT ``AS IS'' AND ANY
-- EXPRESS OR IMPLIED WARRANTIES, INCLUDING, BUT NOT LIMITED TO,
-- THE IMPLIED WARRANTIES OF MERCHANTABILITY AND FITNESS FOR A
-- PARTICULAR PURPOSE ARE DISCLAIMED. IN NO EVENT SHALL THE
-- ZPU PROJECT OR CONTRIBUTORS BE LIABLE FOR ANY DIRECT,
-- INDIRECT, INCIDENTAL, SPECIAL, EXEMPLARY, OR CONSEQUENTIAL DAMAGES
-- (INCLUDING, BUT NOT LIMITED TO, PROCUREMENT OF SUBSTITUTE GOODS
-- OR SERVICES; LOSS OF USE, DATA, OR PROFITS; OR BUSINESS INTERRUPTION)
-- HOWEVER CAUSED AND ON ANY THEORY OF LIABILITY, WHETHER IN CONTRACT,
-- STRICT LIABILITY, OR TORT (INCLUDING NEGLIGENCE OR OTHERWISE)
-- ARISING IN ANY WAY OUT OF THE USE OF THIS SOFTWARE, EVEN IF
-- ADVISED OF THE POSSIBILITY OF SUCH DAMAGE.
-- 
-- The views and conclusions contained in the software and documentation
-- are those of the authors and should not be interpreted as representing
-- official policies, either expressed or implied, of the ZPU Project.

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;


library work;
use work.zpu_config.all;
use work.zpupkg.all;

entity SDBootstrap_ROM is
generic
	(
		maxAddrBitBRAM : integer := maxAddrBitBRAMLimit -- Specify your actual ROM size to save LEs and unnecessary block RAM usage.
	);
port (
	clk : in std_logic;
	areset : in std_logic := '0';
	from_zpu : in ZPU_ToROM;
	to_zpu : out ZPU_FromROM
);
end SDBootstrap_ROM;

architecture arch of SDBootstrap_ROM is

type ram_type is array(natural range 0 to ((2**(maxAddrBitBRAM+1))/4)-1) of std_logic_vector(wordSize-1 downto 0);

shared variable ram : ram_type :=
(
     0 => x"84808080",
     1 => x"ed040000",
     2 => x"00000000",
     3 => x"84808080",
     4 => x"880d8004",
     5 => x"84808080",
     6 => x"940471fd",
     7 => x"06087283",
     8 => x"06098105",
     9 => x"8205832b",
    10 => x"2a83ffff",
    11 => x"06520471",
    12 => x"fc060872",
    13 => x"83060981",
    14 => x"05830510",
    15 => x"10102a81",
    16 => x"ff065204",
    17 => x"71fc0608",
    18 => x"8480809f",
    19 => x"d4738306",
    20 => x"10100508",
    21 => x"067381ff",
    22 => x"06738306",
    23 => x"09810583",
    24 => x"05101010",
    25 => x"2b0772fc",
    26 => x"060c5151",
    27 => x"04028405",
    28 => x"84808080",
    29 => x"880c8480",
    30 => x"8080940b",
    31 => x"8480808d",
    32 => x"8a040000",
    33 => x"02c4050d",
    34 => x"0280c005",
    35 => x"83ffe0e0",
    36 => x"5b568076",
    37 => x"70840558",
    38 => x"08715e5e",
    39 => x"577c7084",
    40 => x"055e0858",
    41 => x"805b7798",
    42 => x"2a78882b",
    43 => x"59547389",
    44 => x"38765e84",
    45 => x"808083d0",
    46 => x"047b802e",
    47 => x"81ea3880",
    48 => x"5c7380e4",
    49 => x"2ea13873",
    50 => x"80e4268e",
    51 => x"387380e3",
    52 => x"2e818738",
    53 => x"84808082",
    54 => x"e8047380",
    55 => x"f32e80e2",
    56 => x"38848080",
    57 => x"82e80475",
    58 => x"84177108",
    59 => x"7e5c5557",
    60 => x"52728025",
    61 => x"8e38ad51",
    62 => x"84808083",
    63 => x"db2d7209",
    64 => x"81055387",
    65 => x"55729c2a",
    66 => x"73842b54",
    67 => x"5271802e",
    68 => x"83388159",
    69 => x"8972258a",
    70 => x"38b71252",
    71 => x"84808082",
    72 => x"a504b012",
    73 => x"5278802e",
    74 => x"89387151",
    75 => x"84808083",
    76 => x"db2dff15",
    77 => x"55748025",
    78 => x"cc388053",
    79 => x"84808083",
    80 => x"81047584",
    81 => x"17710870",
    82 => x"545c5752",
    83 => x"84808083",
    84 => x"ff2d7b53",
    85 => x"84808083",
    86 => x"81047584",
    87 => x"17710856",
    88 => x"57528480",
    89 => x"8083b804",
    90 => x"a5518480",
    91 => x"8083db2d",
    92 => x"73518480",
    93 => x"8083db2d",
    94 => x"82175784",
    95 => x"808083c3",
    96 => x"0472ff14",
    97 => x"54528072",
    98 => x"25b93879",
    99 => x"7081055b",
   100 => x"84808080",
   101 => x"af2d7052",
   102 => x"54848080",
   103 => x"83db2d81",
   104 => x"17578480",
   105 => x"80838104",
   106 => x"73a52e09",
   107 => x"81068938",
   108 => x"815c8480",
   109 => x"8083c304",
   110 => x"73518480",
   111 => x"8083db2d",
   112 => x"81175781",
   113 => x"1b5b837b",
   114 => x"25fddb38",
   115 => x"73fdce38",
   116 => x"7d83ffe0",
   117 => x"800c02bc",
   118 => x"050d0402",
   119 => x"f8050d73",
   120 => x"52c00870",
   121 => x"882a7081",
   122 => x"06515151",
   123 => x"70802ef1",
   124 => x"3871c00c",
   125 => x"7183ffe0",
   126 => x"800c0288",
   127 => x"050d0402",
   128 => x"e8050d80",
   129 => x"78575575",
   130 => x"70840557",
   131 => x"08538054",
   132 => x"72982a73",
   133 => x"882b5452",
   134 => x"71802ea2",
   135 => x"38c00870",
   136 => x"882a7081",
   137 => x"06515151",
   138 => x"70802ef1",
   139 => x"3871c00c",
   140 => x"81158115",
   141 => x"55558374",
   142 => x"25d63871",
   143 => x"ca387483",
   144 => x"ffe0800c",
   145 => x"0298050d",
   146 => x"0402f405",
   147 => x"0d747671",
   148 => x"81ff06d4",
   149 => x"0c535383",
   150 => x"fff1a008",
   151 => x"85387189",
   152 => x"2b527198",
   153 => x"2ad40c71",
   154 => x"902a7081",
   155 => x"ff06d40c",
   156 => x"5171882a",
   157 => x"7081ff06",
   158 => x"d40c5171",
   159 => x"81ff06d4",
   160 => x"0c72902a",
   161 => x"7081ff06",
   162 => x"d40c51d4",
   163 => x"087081ff",
   164 => x"06515182",
   165 => x"b8bf5270",
   166 => x"81ff2e09",
   167 => x"81069438",
   168 => x"81ff0bd4",
   169 => x"0cd40870",
   170 => x"81ff06ff",
   171 => x"14545151",
   172 => x"71e53870",
   173 => x"83ffe080",
   174 => x"0c028c05",
   175 => x"0d0402fc",
   176 => x"050d81c7",
   177 => x"5181ff0b",
   178 => x"d40cff11",
   179 => x"51708025",
   180 => x"f4380284",
   181 => x"050d0402",
   182 => x"f0050d84",
   183 => x"808085be",
   184 => x"2d819c9f",
   185 => x"53805287",
   186 => x"fc80f751",
   187 => x"84808084",
   188 => x"c92d83ff",
   189 => x"e0800854",
   190 => x"83ffe080",
   191 => x"08812e09",
   192 => x"8106ae38",
   193 => x"81ff0bd4",
   194 => x"0c820a52",
   195 => x"849c80e9",
   196 => x"51848080",
   197 => x"84c92d83",
   198 => x"ffe08008",
   199 => x"8e3881ff",
   200 => x"0bd40c73",
   201 => x"53848080",
   202 => x"86b80484",
   203 => x"808085be",
   204 => x"2dff1353",
   205 => x"72ffae38",
   206 => x"7283ffe0",
   207 => x"800c0290",
   208 => x"050d0402",
   209 => x"f4050d81",
   210 => x"ff0bd40c",
   211 => x"8480809f",
   212 => x"e4518480",
   213 => x"8083ff2d",
   214 => x"93538052",
   215 => x"87fc80c1",
   216 => x"51848080",
   217 => x"84c92d83",
   218 => x"ffe08008",
   219 => x"8e3881ff",
   220 => x"0bd40c81",
   221 => x"53848080",
   222 => x"87870484",
   223 => x"808085be",
   224 => x"2dff1353",
   225 => x"72d43872",
   226 => x"83ffe080",
   227 => x"0c028c05",
   228 => x"0d0402f0",
   229 => x"050d8480",
   230 => x"8085be2d",
   231 => x"83aa5284",
   232 => x"9c80c851",
   233 => x"84808084",
   234 => x"c92d83ff",
   235 => x"e0800883",
   236 => x"ffe08008",
   237 => x"53848080",
   238 => x"9ff05254",
   239 => x"84808081",
   240 => x"842d7381",
   241 => x"2e098106",
   242 => x"9038d808",
   243 => x"7083ffff",
   244 => x"06545472",
   245 => x"83aa2ea9",
   246 => x"38848080",
   247 => x"86c32d84",
   248 => x"808087f9",
   249 => x"04815484",
   250 => x"808089b0",
   251 => x"04848080",
   252 => x"a0885184",
   253 => x"80808184",
   254 => x"2d805484",
   255 => x"808089b0",
   256 => x"04735284",
   257 => x"8080a0a4",
   258 => x"51848080",
   259 => x"81842d81",
   260 => x"ff0bd40c",
   261 => x"b1538480",
   262 => x"8085d72d",
   263 => x"83ffe080",
   264 => x"08802e80",
   265 => x"fc388052",
   266 => x"87fc80fa",
   267 => x"51848080",
   268 => x"84c92d83",
   269 => x"ffe08008",
   270 => x"80d53883",
   271 => x"ffe08008",
   272 => x"52848080",
   273 => x"a0bc5184",
   274 => x"80808184",
   275 => x"2d81ff0b",
   276 => x"d40cd408",
   277 => x"81ff0670",
   278 => x"53848080",
   279 => x"a0c85254",
   280 => x"84808081",
   281 => x"842d81ff",
   282 => x"0bd40c81",
   283 => x"ff0bd40c",
   284 => x"81ff0bd4",
   285 => x"0c81ff0b",
   286 => x"d40c7386",
   287 => x"2a708106",
   288 => x"70565153",
   289 => x"72802ea8",
   290 => x"38848080",
   291 => x"87e50483",
   292 => x"ffe08008",
   293 => x"52848080",
   294 => x"a0bc5184",
   295 => x"80808184",
   296 => x"2d72822e",
   297 => x"fec738ff",
   298 => x"135372fe",
   299 => x"e9387254",
   300 => x"7383ffe0",
   301 => x"800c0290",
   302 => x"050d0402",
   303 => x"f4050d81",
   304 => x"0b83fff1",
   305 => x"a00cd008",
   306 => x"708f2a70",
   307 => x"81065151",
   308 => x"5372f338",
   309 => x"72d00c84",
   310 => x"808085be",
   311 => x"2dd00870",
   312 => x"8f2a7081",
   313 => x"06515153",
   314 => x"72f33881",
   315 => x"0bd00c87",
   316 => x"53805284",
   317 => x"d480c051",
   318 => x"84808084",
   319 => x"c92d83ff",
   320 => x"e0800881",
   321 => x"2e973872",
   322 => x"822e0981",
   323 => x"06893880",
   324 => x"53848080",
   325 => x"8ad704ff",
   326 => x"135372d5",
   327 => x"38848080",
   328 => x"87922d83",
   329 => x"ffe08008",
   330 => x"83fff1a0",
   331 => x"0c815287",
   332 => x"fc80d051",
   333 => x"84808084",
   334 => x"c92d81ff",
   335 => x"0bd40cd0",
   336 => x"08708f2a",
   337 => x"70810651",
   338 => x"515372f3",
   339 => x"3872d00c",
   340 => x"81ff0bd4",
   341 => x"0c815372",
   342 => x"83ffe080",
   343 => x"0c028c05",
   344 => x"0d04800b",
   345 => x"83ffe080",
   346 => x"0c0402e0",
   347 => x"050d797b",
   348 => x"57578058",
   349 => x"81ff0bd4",
   350 => x"0cd00870",
   351 => x"8f2a7081",
   352 => x"06515154",
   353 => x"73f33882",
   354 => x"810bd00c",
   355 => x"81ff0bd4",
   356 => x"0c765287",
   357 => x"fc80d151",
   358 => x"84808084",
   359 => x"c92d80db",
   360 => x"c6df5583",
   361 => x"ffe08008",
   362 => x"802e9b38",
   363 => x"83ffe080",
   364 => x"08537652",
   365 => x"848080a0",
   366 => x"d8518480",
   367 => x"8081842d",
   368 => x"8480808c",
   369 => x"930481ff",
   370 => x"0bd40cd4",
   371 => x"087081ff",
   372 => x"06515473",
   373 => x"81fe2e09",
   374 => x"81069c38",
   375 => x"80ff55d8",
   376 => x"08767084",
   377 => x"05580cff",
   378 => x"15557480",
   379 => x"25f13881",
   380 => x"58848080",
   381 => x"8bfd04ff",
   382 => x"155574ca",
   383 => x"3881ff0b",
   384 => x"d40cd008",
   385 => x"708f2a70",
   386 => x"81065151",
   387 => x"5473f338",
   388 => x"73d00c77",
   389 => x"83ffe080",
   390 => x"0c02a005",
   391 => x"0d0402f4",
   392 => x"050d7470",
   393 => x"882a83fe",
   394 => x"80067072",
   395 => x"982a0772",
   396 => x"882b87fc",
   397 => x"80800673",
   398 => x"982b81f0",
   399 => x"0a067173",
   400 => x"070783ff",
   401 => x"e0800c56",
   402 => x"51535102",
   403 => x"8c050d04",
   404 => x"02f8050d",
   405 => x"028e0584",
   406 => x"808080af",
   407 => x"2d74982b",
   408 => x"71902b07",
   409 => x"70902c83",
   410 => x"ffe0800c",
   411 => x"52520288",
   412 => x"050d0402",
   413 => x"f8050d73",
   414 => x"70902b71",
   415 => x"902a0783",
   416 => x"ffe0800c",
   417 => x"52028805",
   418 => x"0d0402ec",
   419 => x"050d800b",
   420 => x"fc800c84",
   421 => x"8080a0f8",
   422 => x"51848080",
   423 => x"83ff2d84",
   424 => x"808089bb",
   425 => x"2d83ffe0",
   426 => x"8008802e",
   427 => x"81f73884",
   428 => x"8080a190",
   429 => x"51848080",
   430 => x"83ff2d84",
   431 => x"80809089",
   432 => x"2d83ffe1",
   433 => x"a0528480",
   434 => x"80a1a851",
   435 => x"8480809c",
   436 => x"ec2d83ff",
   437 => x"e0800880",
   438 => x"2e81ca38",
   439 => x"83ffe1a0",
   440 => x"0b848080",
   441 => x"a1b45254",
   442 => x"84808083",
   443 => x"ff2d8055",
   444 => x"73708105",
   445 => x"55848080",
   446 => x"80af2d53",
   447 => x"72a02e80",
   448 => x"e33872a3",
   449 => x"2e818438",
   450 => x"7280c72e",
   451 => x"0981068d",
   452 => x"38848080",
   453 => x"808c2d84",
   454 => x"80808ebf",
   455 => x"04728a2e",
   456 => x"0981068d",
   457 => x"38848080",
   458 => x"80942d84",
   459 => x"80808ebf",
   460 => x"047280cc",
   461 => x"2e098106",
   462 => x"863883ff",
   463 => x"e1a05472",
   464 => x"81df06f0",
   465 => x"057081ff",
   466 => x"065153b8",
   467 => x"73278938",
   468 => x"ef137081",
   469 => x"ff065153",
   470 => x"74842b73",
   471 => x"07558480",
   472 => x"808df004",
   473 => x"72a32ea3",
   474 => x"38737081",
   475 => x"05558480",
   476 => x"8080af2d",
   477 => x"5372a02e",
   478 => x"f038ff14",
   479 => x"75537052",
   480 => x"54848080",
   481 => x"9cec2d74",
   482 => x"fc800c73",
   483 => x"70810555",
   484 => x"84808080",
   485 => x"af2d5372",
   486 => x"8a2e0981",
   487 => x"06ed3884",
   488 => x"80808dee",
   489 => x"04848080",
   490 => x"a1c85184",
   491 => x"808083ff",
   492 => x"2d800b83",
   493 => x"ffe0800c",
   494 => x"0294050d",
   495 => x"0402e805",
   496 => x"0d77797b",
   497 => x"58555580",
   498 => x"53727625",
   499 => x"af387470",
   500 => x"81055684",
   501 => x"808080af",
   502 => x"2d747081",
   503 => x"05568480",
   504 => x"8080af2d",
   505 => x"52527171",
   506 => x"2e893881",
   507 => x"51848080",
   508 => x"8ffe0481",
   509 => x"13538480",
   510 => x"808fc904",
   511 => x"80517083",
   512 => x"ffe0800c",
   513 => x"0298050d",
   514 => x"0402d805",
   515 => x"0dff0b83",
   516 => x"fff5cc0c",
   517 => x"800b83ff",
   518 => x"f5e00c84",
   519 => x"8080a1d4",
   520 => x"51848080",
   521 => x"83ff2d83",
   522 => x"fff1b852",
   523 => x"80518480",
   524 => x"808aea2d",
   525 => x"83ffe080",
   526 => x"085483ff",
   527 => x"e0800895",
   528 => x"38848080",
   529 => x"a1e45184",
   530 => x"808083ff",
   531 => x"2d735584",
   532 => x"808098ae",
   533 => x"04848080",
   534 => x"a1f85184",
   535 => x"808083ff",
   536 => x"2d805681",
   537 => x"0b83fff1",
   538 => x"ac0c8853",
   539 => x"848080a2",
   540 => x"905283ff",
   541 => x"f1ee5184",
   542 => x"80808fbd",
   543 => x"2d83ffe0",
   544 => x"8008762e",
   545 => x"0981068b",
   546 => x"3883ffe0",
   547 => x"800883ff",
   548 => x"f1ac0c88",
   549 => x"53848080",
   550 => x"a29c5283",
   551 => x"fff28a51",
   552 => x"8480808f",
   553 => x"bd2d83ff",
   554 => x"e080088b",
   555 => x"3883ffe0",
   556 => x"800883ff",
   557 => x"f1ac0c83",
   558 => x"fff1ac08",
   559 => x"52848080",
   560 => x"a2a85184",
   561 => x"80808184",
   562 => x"2d83fff1",
   563 => x"ac08802e",
   564 => x"81cb3883",
   565 => x"fff4fe0b",
   566 => x"84808080",
   567 => x"af2d83ff",
   568 => x"f4ff0b84",
   569 => x"808080af",
   570 => x"2d71982b",
   571 => x"71902b07",
   572 => x"83fff580",
   573 => x"0b848080",
   574 => x"80af2d70",
   575 => x"882b7207",
   576 => x"83fff581",
   577 => x"0b848080",
   578 => x"80af2d71",
   579 => x"0783fff5",
   580 => x"b60b8480",
   581 => x"8080af2d",
   582 => x"83fff5b7",
   583 => x"0b848080",
   584 => x"80af2d71",
   585 => x"882b0753",
   586 => x"5f54525a",
   587 => x"56575573",
   588 => x"81abaa2e",
   589 => x"09810695",
   590 => x"38755184",
   591 => x"80808c9e",
   592 => x"2d83ffe0",
   593 => x"80085684",
   594 => x"808092e6",
   595 => x"047382d4",
   596 => x"d52e9338",
   597 => x"848080a2",
   598 => x"bc518480",
   599 => x"8083ff2d",
   600 => x"84808094",
   601 => x"f2047552",
   602 => x"848080a2",
   603 => x"dc518480",
   604 => x"8081842d",
   605 => x"83fff1b8",
   606 => x"52755184",
   607 => x"80808aea",
   608 => x"2d83ffe0",
   609 => x"80085583",
   610 => x"ffe08008",
   611 => x"802e859e",
   612 => x"38848080",
   613 => x"a2f45184",
   614 => x"808083ff",
   615 => x"2d848080",
   616 => x"a39c5184",
   617 => x"80808184",
   618 => x"2d885384",
   619 => x"8080a29c",
   620 => x"5283fff2",
   621 => x"8a518480",
   622 => x"808fbd2d",
   623 => x"83ffe080",
   624 => x"088e3881",
   625 => x"0b83fff5",
   626 => x"e00c8480",
   627 => x"8093fe04",
   628 => x"88538480",
   629 => x"80a29052",
   630 => x"83fff1ee",
   631 => x"51848080",
   632 => x"8fbd2d83",
   633 => x"ffe08008",
   634 => x"802e9338",
   635 => x"848080a3",
   636 => x"b4518480",
   637 => x"8081842d",
   638 => x"84808094",
   639 => x"f20483ff",
   640 => x"f5b60b84",
   641 => x"808080af",
   642 => x"2d547380",
   643 => x"d52e0981",
   644 => x"0680df38",
   645 => x"83fff5b7",
   646 => x"0b848080",
   647 => x"80af2d54",
   648 => x"7381aa2e",
   649 => x"09810680",
   650 => x"c938800b",
   651 => x"83fff1b8",
   652 => x"0b848080",
   653 => x"80af2d56",
   654 => x"547481e9",
   655 => x"2e833881",
   656 => x"547481eb",
   657 => x"2e8c3880",
   658 => x"5573752e",
   659 => x"09810683",
   660 => x"dd3883ff",
   661 => x"f1c30b84",
   662 => x"808080af",
   663 => x"2d557492",
   664 => x"3883fff1",
   665 => x"c40b8480",
   666 => x"8080af2d",
   667 => x"5473822e",
   668 => x"89388055",
   669 => x"84808098",
   670 => x"ae0483ff",
   671 => x"f1c50b84",
   672 => x"808080af",
   673 => x"2d7083ff",
   674 => x"f5e80cff",
   675 => x"0583fff5",
   676 => x"dc0c83ff",
   677 => x"f1c60b84",
   678 => x"808080af",
   679 => x"2d83fff1",
   680 => x"c70b8480",
   681 => x"8080af2d",
   682 => x"58760577",
   683 => x"82802905",
   684 => x"7083fff5",
   685 => x"d00c83ff",
   686 => x"f1c80b84",
   687 => x"808080af",
   688 => x"2d7083ff",
   689 => x"f5c80c83",
   690 => x"fff5e008",
   691 => x"59575876",
   692 => x"802e81ea",
   693 => x"38885384",
   694 => x"8080a29c",
   695 => x"5283fff2",
   696 => x"8a518480",
   697 => x"808fbd2d",
   698 => x"83ffe080",
   699 => x"0882bf38",
   700 => x"83fff5e8",
   701 => x"0870842b",
   702 => x"83fff5b8",
   703 => x"0c7083ff",
   704 => x"f5e40c83",
   705 => x"fff1dd0b",
   706 => x"84808080",
   707 => x"af2d83ff",
   708 => x"f1dc0b84",
   709 => x"808080af",
   710 => x"2d718280",
   711 => x"290583ff",
   712 => x"f1de0b84",
   713 => x"808080af",
   714 => x"2d708480",
   715 => x"80291283",
   716 => x"fff1df0b",
   717 => x"84808080",
   718 => x"af2d7081",
   719 => x"800a2912",
   720 => x"7083fff1",
   721 => x"b00c83ff",
   722 => x"f5c80871",
   723 => x"2983fff5",
   724 => x"d0080570",
   725 => x"83fff5f0",
   726 => x"0c83fff1",
   727 => x"e50b8480",
   728 => x"8080af2d",
   729 => x"83fff1e4",
   730 => x"0b848080",
   731 => x"80af2d71",
   732 => x"82802905",
   733 => x"83fff1e6",
   734 => x"0b848080",
   735 => x"80af2d70",
   736 => x"84808029",
   737 => x"1283fff1",
   738 => x"e70b8480",
   739 => x"8080af2d",
   740 => x"70982b81",
   741 => x"f00a0672",
   742 => x"057083ff",
   743 => x"f1b40cfe",
   744 => x"117e2977",
   745 => x"0583fff5",
   746 => x"d80c5259",
   747 => x"5243545e",
   748 => x"51525952",
   749 => x"5d575957",
   750 => x"84808098",
   751 => x"ac0483ff",
   752 => x"f1ca0b84",
   753 => x"808080af",
   754 => x"2d83fff1",
   755 => x"c90b8480",
   756 => x"8080af2d",
   757 => x"71828029",
   758 => x"057083ff",
   759 => x"f5b80c70",
   760 => x"a02983ff",
   761 => x"0570892a",
   762 => x"7083fff5",
   763 => x"e40c83ff",
   764 => x"f1cf0b84",
   765 => x"808080af",
   766 => x"2d83fff1",
   767 => x"ce0b8480",
   768 => x"8080af2d",
   769 => x"71828029",
   770 => x"057083ff",
   771 => x"f1b00c7b",
   772 => x"71291e70",
   773 => x"83fff5d8",
   774 => x"0c7d83ff",
   775 => x"f1b40c73",
   776 => x"0583fff5",
   777 => x"f00c555e",
   778 => x"51515555",
   779 => x"81557483",
   780 => x"ffe0800c",
   781 => x"02a8050d",
   782 => x"0402ec05",
   783 => x"0d767087",
   784 => x"2c7180ff",
   785 => x"06575553",
   786 => x"83fff5e0",
   787 => x"088a3872",
   788 => x"882c7381",
   789 => x"ff065654",
   790 => x"7383fff5",
   791 => x"cc082ea9",
   792 => x"3883fff1",
   793 => x"b85283ff",
   794 => x"f5d00814",
   795 => x"51848080",
   796 => x"8aea2d83",
   797 => x"ffe08008",
   798 => x"5383ffe0",
   799 => x"8008802e",
   800 => x"80cf3873",
   801 => x"83fff5cc",
   802 => x"0c83fff5",
   803 => x"e008802e",
   804 => x"a2387484",
   805 => x"2983fff1",
   806 => x"b8057008",
   807 => x"52538480",
   808 => x"808c9e2d",
   809 => x"83ffe080",
   810 => x"08f00a06",
   811 => x"55848080",
   812 => x"99cf0474",
   813 => x"1083fff1",
   814 => x"b8057084",
   815 => x"8080809a",
   816 => x"2d525384",
   817 => x"80808cd0",
   818 => x"2d83ffe0",
   819 => x"80085574",
   820 => x"537283ff",
   821 => x"e0800c02",
   822 => x"94050d04",
   823 => x"02cc050d",
   824 => x"7e605e5b",
   825 => x"8056ff0b",
   826 => x"83fff5cc",
   827 => x"0c83fff1",
   828 => x"b40883ff",
   829 => x"f5d80856",
   830 => x"5783fff5",
   831 => x"e008762e",
   832 => x"8f3883ff",
   833 => x"f5e80884",
   834 => x"2b598480",
   835 => x"809a9804",
   836 => x"83fff5e4",
   837 => x"08842b59",
   838 => x"805a7979",
   839 => x"2781f038",
   840 => x"798f06a0",
   841 => x"17575473",
   842 => x"a4387452",
   843 => x"848080a3",
   844 => x"d4518480",
   845 => x"8081842d",
   846 => x"83fff1b8",
   847 => x"52745181",
   848 => x"15558480",
   849 => x"808aea2d",
   850 => x"83fff1b8",
   851 => x"56807684",
   852 => x"808080af",
   853 => x"2d555873",
   854 => x"782e8338",
   855 => x"81587381",
   856 => x"e52e81a2",
   857 => x"38817079",
   858 => x"06555c73",
   859 => x"802e8196",
   860 => x"388b1684",
   861 => x"808080af",
   862 => x"2d980658",
   863 => x"77818738",
   864 => x"8b537c52",
   865 => x"75518480",
   866 => x"808fbd2d",
   867 => x"83ffe080",
   868 => x"0880f338",
   869 => x"9c160851",
   870 => x"8480808c",
   871 => x"9e2d83ff",
   872 => x"e0800884",
   873 => x"1c0c9a16",
   874 => x"84808080",
   875 => x"9a2d5184",
   876 => x"80808cd0",
   877 => x"2d83ffe0",
   878 => x"800883ff",
   879 => x"e0800855",
   880 => x"5583fff5",
   881 => x"e008802e",
   882 => x"a0389416",
   883 => x"84808080",
   884 => x"9a2d5184",
   885 => x"80808cd0",
   886 => x"2d83ffe0",
   887 => x"8008902b",
   888 => x"83fff00a",
   889 => x"06701651",
   890 => x"5473881c",
   891 => x"0c777b0c",
   892 => x"7c528480",
   893 => x"80a3f451",
   894 => x"84808081",
   895 => x"842d7b54",
   896 => x"8480809c",
   897 => x"e104811a",
   898 => x"5a848080",
   899 => x"9a9a0483",
   900 => x"fff5e008",
   901 => x"802e80c7",
   902 => x"38765184",
   903 => x"808098b9",
   904 => x"2d83ffe0",
   905 => x"800883ff",
   906 => x"e0800853",
   907 => x"848080a4",
   908 => x"88525784",
   909 => x"80808184",
   910 => x"2d7680ff",
   911 => x"fffff806",
   912 => x"547380ff",
   913 => x"fffff82e",
   914 => x"9638fe17",
   915 => x"83fff5e8",
   916 => x"082983ff",
   917 => x"f5f00805",
   918 => x"55848080",
   919 => x"9a980480",
   920 => x"547383ff",
   921 => x"e0800c02",
   922 => x"b4050d04",
   923 => x"02e4050d",
   924 => x"787a7154",
   925 => x"83fff5bc",
   926 => x"53555584",
   927 => x"808099dc",
   928 => x"2d83ffe0",
   929 => x"800881ff",
   930 => x"06537280",
   931 => x"2e818838",
   932 => x"848080a4",
   933 => x"a0518480",
   934 => x"8083ff2d",
   935 => x"83fff5c0",
   936 => x"0883ff05",
   937 => x"892a5780",
   938 => x"70565675",
   939 => x"77258187",
   940 => x"3883fff5",
   941 => x"c408fe05",
   942 => x"83fff5e8",
   943 => x"082983ff",
   944 => x"f5f00811",
   945 => x"7683fff5",
   946 => x"dc080605",
   947 => x"75545253",
   948 => x"8480808a",
   949 => x"ea2d83ff",
   950 => x"e0800880",
   951 => x"2e80cc38",
   952 => x"81157083",
   953 => x"fff5dc08",
   954 => x"06545572",
   955 => x"973883ff",
   956 => x"f5c40851",
   957 => x"84808098",
   958 => x"b92d83ff",
   959 => x"e0800883",
   960 => x"fff5c40c",
   961 => x"84801481",
   962 => x"17575476",
   963 => x"7624ffa1",
   964 => x"38848080",
   965 => x"9eb70474",
   966 => x"52848080",
   967 => x"a4bc5184",
   968 => x"80808184",
   969 => x"2d848080",
   970 => x"9eb90483",
   971 => x"ffe08008",
   972 => x"53848080",
   973 => x"9eb90481",
   974 => x"537283ff",
   975 => x"e0800c02",
   976 => x"9c050d04",
   977 => x"83ffe08c",
   978 => x"080283ff",
   979 => x"e08c0cff",
   980 => x"3d0d800b",
   981 => x"83ffe08c",
   982 => x"08fc050c",
   983 => x"83ffe08c",
   984 => x"08880508",
   985 => x"8106ff11",
   986 => x"70097083",
   987 => x"ffe08c08",
   988 => x"8c050806",
   989 => x"83ffe08c",
   990 => x"08fc0508",
   991 => x"1183ffe0",
   992 => x"8c08fc05",
   993 => x"0c83ffe0",
   994 => x"8c088805",
   995 => x"08812a83",
   996 => x"ffe08c08",
   997 => x"88050c83",
   998 => x"ffe08c08",
   999 => x"8c050810",
  1000 => x"83ffe08c",
  1001 => x"088c050c",
  1002 => x"51515151",
  1003 => x"83ffe08c",
  1004 => x"08880508",
  1005 => x"802e8438",
  1006 => x"ffa23983",
  1007 => x"ffe08c08",
  1008 => x"fc050870",
  1009 => x"83ffe080",
  1010 => x"0c51833d",
  1011 => x"0d83ffe0",
  1012 => x"8c0c0400",
  1013 => x"00ffffff",
  1014 => x"ff00ffff",
  1015 => x"ffff00ff",
  1016 => x"ffffff00",
  1017 => x"436d645f",
  1018 => x"696e6974",
  1019 => x"0a000000",
  1020 => x"636d645f",
  1021 => x"434d4438",
  1022 => x"20726573",
  1023 => x"706f6e73",
  1024 => x"653a2025",
  1025 => x"640a0000",
  1026 => x"53444843",
  1027 => x"20496e69",
  1028 => x"7469616c",
  1029 => x"697a6174",
  1030 => x"696f6e20",
  1031 => x"6572726f",
  1032 => x"72210a00",
  1033 => x"434d4438",
  1034 => x"5f342072",
  1035 => x"6573706f",
  1036 => x"6e73653a",
  1037 => x"2025640a",
  1038 => x"00000000",
  1039 => x"434d4435",
  1040 => x"38202564",
  1041 => x"0a202000",
  1042 => x"434d4435",
  1043 => x"385f3220",
  1044 => x"25640a20",
  1045 => x"20000000",
  1046 => x"52656164",
  1047 => x"20636f6d",
  1048 => x"6d616e64",
  1049 => x"20666169",
  1050 => x"6c656420",
  1051 => x"61742025",
  1052 => x"64202825",
  1053 => x"64290a00",
  1054 => x"496e6974",
  1055 => x"69616c69",
  1056 => x"7a696e67",
  1057 => x"20534420",
  1058 => x"63617264",
  1059 => x"0a000000",
  1060 => x"48756e74",
  1061 => x"696e6720",
  1062 => x"666f7220",
  1063 => x"70617274",
  1064 => x"6974696f",
  1065 => x"6e0a0000",
  1066 => x"4d414e49",
  1067 => x"46455354",
  1068 => x"4d535400",
  1069 => x"50617273",
  1070 => x"696e6720",
  1071 => x"6d616e69",
  1072 => x"66657374",
  1073 => x"0a000000",
  1074 => x"52657475",
  1075 => x"726e696e",
  1076 => x"670a0000",
  1077 => x"52656164",
  1078 => x"696e6720",
  1079 => x"4d42520a",
  1080 => x"00000000",
  1081 => x"52656164",
  1082 => x"206f6620",
  1083 => x"4d425220",
  1084 => x"6661696c",
  1085 => x"65640a00",
  1086 => x"4d425220",
  1087 => x"73756363",
  1088 => x"65737366",
  1089 => x"756c6c79",
  1090 => x"20726561",
  1091 => x"640a0000",
  1092 => x"46415431",
  1093 => x"36202020",
  1094 => x"00000000",
  1095 => x"46415433",
  1096 => x"32202020",
  1097 => x"00000000",
  1098 => x"50617274",
  1099 => x"6974696f",
  1100 => x"6e636f75",
  1101 => x"6e742025",
  1102 => x"640a0000",
  1103 => x"4e6f2070",
  1104 => x"61727469",
  1105 => x"74696f6e",
  1106 => x"20736967",
  1107 => x"6e617475",
  1108 => x"72652066",
  1109 => x"6f756e64",
  1110 => x"0a000000",
  1111 => x"52656164",
  1112 => x"696e6720",
  1113 => x"626f6f74",
  1114 => x"20736563",
  1115 => x"746f7220",
  1116 => x"25640a00",
  1117 => x"52656164",
  1118 => x"20626f6f",
  1119 => x"74207365",
  1120 => x"63746f72",
  1121 => x"2066726f",
  1122 => x"6d206669",
  1123 => x"72737420",
  1124 => x"70617274",
  1125 => x"6974696f",
  1126 => x"6e0a0000",
  1127 => x"48756e74",
  1128 => x"696e6720",
  1129 => x"666f7220",
  1130 => x"66696c65",
  1131 => x"73797374",
  1132 => x"656d0a00",
  1133 => x"556e7375",
  1134 => x"70706f72",
  1135 => x"74656420",
  1136 => x"70617274",
  1137 => x"6974696f",
  1138 => x"6e207479",
  1139 => x"7065210d",
  1140 => x"00000000",
  1141 => x"52656164",
  1142 => x"696e6720",
  1143 => x"64697265",
  1144 => x"63746f72",
  1145 => x"79207365",
  1146 => x"63746f72",
  1147 => x"2025640a",
  1148 => x"00000000",
  1149 => x"66696c65",
  1150 => x"20222573",
  1151 => x"2220666f",
  1152 => x"756e640d",
  1153 => x"00000000",
  1154 => x"47657446",
  1155 => x"41544c69",
  1156 => x"6e6b2072",
  1157 => x"65747572",
  1158 => x"6e656420",
  1159 => x"25640a00",
  1160 => x"4f70656e",
  1161 => x"65642066",
  1162 => x"696c652c",
  1163 => x"206c6f61",
  1164 => x"64696e67",
  1165 => x"2e2e2e0a",
  1166 => x"00000000",
  1167 => x"43616e27",
  1168 => x"74206f70",
  1169 => x"656e2025",
  1170 => x"730a0000",
	others => x"00000000"
);

begin

process (clk)
begin
	if (clk'event and clk = '1') then
		if (from_zpu.memAWriteEnable = '1') and (from_zpu.memBWriteEnable = '1') and (from_zpu.memAAddr=from_zpu.memBAddr) and (from_zpu.memAWrite/=from_zpu.memBWrite) then
			report "write collision" severity failure;
		end if;
	
		if (from_zpu.memAWriteEnable = '1') then
			ram(to_integer(unsigned(from_zpu.memAAddr(maxAddrBitBRAM downto 2)))) := from_zpu.memAWrite;
			to_zpu.memARead <= from_zpu.memAWrite;
		else
			to_zpu.memARead <= ram(to_integer(unsigned(from_zpu.memAAddr(maxAddrBitBRAM downto 2))));
		end if;
	end if;
end process;

process (clk)
begin
	if (clk'event and clk = '1') then
		if (from_zpu.memBWriteEnable = '1') then
			ram(to_integer(unsigned(from_zpu.memBAddr(maxAddrBitBRAM downto 2)))) := from_zpu.memBWrite;
			to_zpu.memBRead <= from_zpu.memBWrite;
		else
			to_zpu.memBRead <= ram(to_integer(unsigned(from_zpu.memBAddr(maxAddrBitBRAM downto 2))));
		end if;
	end if;
end process;


end arch;

