-- ZPU
--
-- Copyright 2004-2008 oharboe - �yvind Harboe - oyvind.harboe@zylin.com
-- Modified by Alastair M. Robinson for the ZPUFlex project.
--
-- The FreeBSD license
-- 
-- Redistribution and use in source and binary forms, with or without
-- modification, are permitted provided that the following conditions
-- are met:
-- 
-- 1. Redistributions of source code must retain the above copyright
--    notice, this list of conditions and the following disclaimer.
-- 2. Redistributions in binary form must reproduce the above
--    copyright notice, this list of conditions and the following
--    disclaimer in the documentation and/or other materials
--    provided with the distribution.
-- 
-- THIS SOFTWARE IS PROVIDED BY THE ZPU PROJECT ``AS IS'' AND ANY
-- EXPRESS OR IMPLIED WARRANTIES, INCLUDING, BUT NOT LIMITED TO,
-- THE IMPLIED WARRANTIES OF MERCHANTABILITY AND FITNESS FOR A
-- PARTICULAR PURPOSE ARE DISCLAIMED. IN NO EVENT SHALL THE
-- ZPU PROJECT OR CONTRIBUTORS BE LIABLE FOR ANY DIRECT,
-- INDIRECT, INCIDENTAL, SPECIAL, EXEMPLARY, OR CONSEQUENTIAL DAMAGES
-- (INCLUDING, BUT NOT LIMITED TO, PROCUREMENT OF SUBSTITUTE GOODS
-- OR SERVICES; LOSS OF USE, DATA, OR PROFITS; OR BUSINESS INTERRUPTION)
-- HOWEVER CAUSED AND ON ANY THEORY OF LIABILITY, WHETHER IN CONTRACT,
-- STRICT LIABILITY, OR TORT (INCLUDING NEGLIGENCE OR OTHERWISE)
-- ARISING IN ANY WAY OUT OF THE USE OF THIS SOFTWARE, EVEN IF
-- ADVISED OF THE POSSIBILITY OF SUCH DAMAGE.
-- 
-- The views and conclusions contained in the software and documentation
-- are those of the authors and should not be interpreted as representing
-- official policies, either expressed or implied, of the ZPU Project.

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;


library work;
use work.zpu_config.all;
use work.zpupkg.all;

entity VGATest_ROM is
generic
	(
		maxAddrBitBRAM : integer := maxAddrBitBRAMLimit -- Specify your actual ROM size to save LEs and unnecessary block RAM usage.
	);
port (
	clk : in std_logic;
	areset : in std_logic := '0';
	from_zpu : in ZPU_ToROM;
	to_zpu : out ZPU_FromROM
);
end VGATest_ROM;

architecture arch of VGATest_ROM is

type ram_type is array(natural range 0 to ((2**(maxAddrBitBRAM+1))/4)-1) of std_logic_vector(wordSize-1 downto 0);

shared variable ram : ram_type :=
(
     0 => x"0b0b0b88",
     1 => x"dd040000",
     2 => x"00000000",
     3 => x"00000000",
     4 => x"00000000",
     5 => x"00000000",
     6 => x"00000000",
     7 => x"00000000",
     8 => x"88088c08",
     9 => x"90080b0b",
    10 => x"0b88e708",
    11 => x"2d900c8c",
    12 => x"0c880c04",
    13 => x"00000000",
    14 => x"00000000",
    15 => x"00000000",
    16 => x"71fd0608",
    17 => x"72830609",
    18 => x"81058205",
    19 => x"832b2a83",
    20 => x"ffff0652",
    21 => x"04000000",
    22 => x"00000000",
    23 => x"00000000",
    24 => x"71fd0608",
    25 => x"83ffff73",
    26 => x"83060981",
    27 => x"05820583",
    28 => x"2b2b0906",
    29 => x"7383ffff",
    30 => x"0b0b0b0b",
    31 => x"83a50400",
    32 => x"72098105",
    33 => x"72057373",
    34 => x"09060906",
    35 => x"73097306",
    36 => x"070a8106",
    37 => x"53510400",
    38 => x"00000000",
    39 => x"00000000",
    40 => x"72722473",
    41 => x"732e0753",
    42 => x"51040000",
    43 => x"00000000",
    44 => x"00000000",
    45 => x"00000000",
    46 => x"00000000",
    47 => x"00000000",
    48 => x"71737109",
    49 => x"71068106",
    50 => x"09810572",
    51 => x"0a100a72",
    52 => x"0a100a31",
    53 => x"050a8106",
    54 => x"51515351",
    55 => x"04000000",
    56 => x"72722673",
    57 => x"732e0753",
    58 => x"51040000",
    59 => x"00000000",
    60 => x"00000000",
    61 => x"00000000",
    62 => x"00000000",
    63 => x"00000000",
    64 => x"00000000",
    65 => x"00000000",
    66 => x"00000000",
    67 => x"00000000",
    68 => x"00000000",
    69 => x"00000000",
    70 => x"00000000",
    71 => x"00000000",
    72 => x"0b0b0b88",
    73 => x"ba040000",
    74 => x"00000000",
    75 => x"00000000",
    76 => x"00000000",
    77 => x"00000000",
    78 => x"00000000",
    79 => x"00000000",
    80 => x"720a722b",
    81 => x"0a535104",
    82 => x"00000000",
    83 => x"00000000",
    84 => x"00000000",
    85 => x"00000000",
    86 => x"00000000",
    87 => x"00000000",
    88 => x"72729f06",
    89 => x"0981050b",
    90 => x"0b0b889f",
    91 => x"05040000",
    92 => x"00000000",
    93 => x"00000000",
    94 => x"00000000",
    95 => x"00000000",
    96 => x"72722aff",
    97 => x"739f062a",
    98 => x"0974090a",
    99 => x"8106ff05",
   100 => x"06075351",
   101 => x"04000000",
   102 => x"00000000",
   103 => x"00000000",
   104 => x"71715351",
   105 => x"04067383",
   106 => x"06098105",
   107 => x"8205832b",
   108 => x"0b2b0772",
   109 => x"fc060c51",
   110 => x"51040000",
   111 => x"00000000",
   112 => x"72098105",
   113 => x"72050970",
   114 => x"81050906",
   115 => x"0a810653",
   116 => x"51040000",
   117 => x"00000000",
   118 => x"00000000",
   119 => x"00000000",
   120 => x"72098105",
   121 => x"72050970",
   122 => x"81050906",
   123 => x"0a098106",
   124 => x"53510400",
   125 => x"00000000",
   126 => x"00000000",
   127 => x"00000000",
   128 => x"71098105",
   129 => x"52040000",
   130 => x"00000000",
   131 => x"00000000",
   132 => x"00000000",
   133 => x"00000000",
   134 => x"00000000",
   135 => x"00000000",
   136 => x"72720981",
   137 => x"05055351",
   138 => x"04000000",
   139 => x"00000000",
   140 => x"00000000",
   141 => x"00000000",
   142 => x"00000000",
   143 => x"00000000",
   144 => x"72097206",
   145 => x"73730906",
   146 => x"07535104",
   147 => x"00000000",
   148 => x"00000000",
   149 => x"00000000",
   150 => x"00000000",
   151 => x"00000000",
   152 => x"71fc0608",
   153 => x"72830609",
   154 => x"81058305",
   155 => x"1010102a",
   156 => x"81ff0652",
   157 => x"04000000",
   158 => x"00000000",
   159 => x"00000000",
   160 => x"71fc0608",
   161 => x"0b0b0b91",
   162 => x"e4738306",
   163 => x"10100508",
   164 => x"060b0b0b",
   165 => x"88a20400",
   166 => x"00000000",
   167 => x"00000000",
   168 => x"88088c08",
   169 => x"90087575",
   170 => x"0b0b0b8d",
   171 => x"e52d5050",
   172 => x"88085690",
   173 => x"0c8c0c88",
   174 => x"0c510400",
   175 => x"00000000",
   176 => x"88088c08",
   177 => x"90087575",
   178 => x"0b0b0b8f",
   179 => x"972d5050",
   180 => x"88085690",
   181 => x"0c8c0c88",
   182 => x"0c510400",
   183 => x"00000000",
   184 => x"72097081",
   185 => x"0509060a",
   186 => x"8106ff05",
   187 => x"70547106",
   188 => x"73097274",
   189 => x"05ff0506",
   190 => x"07515151",
   191 => x"04000000",
   192 => x"72097081",
   193 => x"0509060a",
   194 => x"098106ff",
   195 => x"05705471",
   196 => x"06730972",
   197 => x"7405ff05",
   198 => x"06075151",
   199 => x"51040000",
   200 => x"05ff0504",
   201 => x"00000000",
   202 => x"00000000",
   203 => x"00000000",
   204 => x"00000000",
   205 => x"00000000",
   206 => x"00000000",
   207 => x"00000000",
   208 => x"04000000",
   209 => x"00000000",
   210 => x"00000000",
   211 => x"00000000",
   212 => x"00000000",
   213 => x"00000000",
   214 => x"00000000",
   215 => x"00000000",
   216 => x"71810552",
   217 => x"04000000",
   218 => x"00000000",
   219 => x"00000000",
   220 => x"00000000",
   221 => x"00000000",
   222 => x"00000000",
   223 => x"00000000",
   224 => x"00000000",
   225 => x"00000000",
   226 => x"00000000",
   227 => x"00000000",
   228 => x"00000000",
   229 => x"00000000",
   230 => x"00000000",
   231 => x"00000000",
   232 => x"02840572",
   233 => x"10100552",
   234 => x"04000000",
   235 => x"00000000",
   236 => x"00000000",
   237 => x"00000000",
   238 => x"00000000",
   239 => x"00000000",
   240 => x"00000000",
   241 => x"00000000",
   242 => x"00000000",
   243 => x"00000000",
   244 => x"00000000",
   245 => x"00000000",
   246 => x"00000000",
   247 => x"00000000",
   248 => x"717105ff",
   249 => x"05715351",
   250 => x"020d0400",
   251 => x"00000000",
   252 => x"00000000",
   253 => x"00000000",
   254 => x"00000000",
   255 => x"00000000",
   256 => x"10101010",
   257 => x"10101010",
   258 => x"10101010",
   259 => x"10101010",
   260 => x"10101010",
   261 => x"10101010",
   262 => x"10101010",
   263 => x"10101053",
   264 => x"51047381",
   265 => x"ff067383",
   266 => x"06098105",
   267 => x"83051010",
   268 => x"102b0772",
   269 => x"fc060c51",
   270 => x"51047272",
   271 => x"80728106",
   272 => x"ff050972",
   273 => x"06057110",
   274 => x"52720a10",
   275 => x"0a5372ed",
   276 => x"38515153",
   277 => x"51040000",
   278 => x"800488da",
   279 => x"0488da0b",
   280 => x"8cd90404",
   281 => x"00000000",
   282 => x"00046302",
   283 => x"c0050d02",
   284 => x"80c4050b",
   285 => x"0b0b92d8",
   286 => x"5a5c807c",
   287 => x"7084055e",
   288 => x"08715f5f",
   289 => x"577d7084",
   290 => x"055f0856",
   291 => x"80587598",
   292 => x"2a76882b",
   293 => x"57557480",
   294 => x"2e82cd38",
   295 => x"7c802eb9",
   296 => x"38805d74",
   297 => x"80e42e81",
   298 => x"9f387480",
   299 => x"e42680dc",
   300 => x"387480e3",
   301 => x"2eba38a5",
   302 => x"518bf12d",
   303 => x"74518bf1",
   304 => x"2d821757",
   305 => x"81185883",
   306 => x"7825c338",
   307 => x"74ffb638",
   308 => x"7e880c02",
   309 => x"80c0050d",
   310 => x"0474a52e",
   311 => x"09810698",
   312 => x"38810b81",
   313 => x"19595d83",
   314 => x"7825ffa2",
   315 => x"3889cc04",
   316 => x"7b841d71",
   317 => x"08575d5a",
   318 => x"74518bf1",
   319 => x"2d811781",
   320 => x"19595783",
   321 => x"7825ff86",
   322 => x"3889cc04",
   323 => x"7480f32e",
   324 => x"098106ff",
   325 => x"a2387b84",
   326 => x"1d710870",
   327 => x"545b5d54",
   328 => x"8c922d80",
   329 => x"0bff1155",
   330 => x"53807325",
   331 => x"ff963878",
   332 => x"7081055a",
   333 => x"84e02d70",
   334 => x"52558bf1",
   335 => x"2d811774",
   336 => x"ff165654",
   337 => x"578aa904",
   338 => x"7b841d71",
   339 => x"080b0b0b",
   340 => x"92d80b0b",
   341 => x"0b0b9288",
   342 => x"615f585e",
   343 => x"525d5372",
   344 => x"ba38b00b",
   345 => x"0b0b0b92",
   346 => x"880b8580",
   347 => x"2d811454",
   348 => x"ff145473",
   349 => x"84e02d7b",
   350 => x"7081055d",
   351 => x"85802d81",
   352 => x"1a5a730b",
   353 => x"0b0b9288",
   354 => x"2e098106",
   355 => x"e338807b",
   356 => x"85802d79",
   357 => x"ff115553",
   358 => x"8aa9048a",
   359 => x"5272518d",
   360 => x"c02d8808",
   361 => x"91f40584",
   362 => x"e02d7470",
   363 => x"81055685",
   364 => x"802d8a52",
   365 => x"72518d9b",
   366 => x"2d880853",
   367 => x"8808dc38",
   368 => x"730b0b0b",
   369 => x"92882ec6",
   370 => x"38ff1454",
   371 => x"7384e02d",
   372 => x"7b708105",
   373 => x"5d85802d",
   374 => x"811a5a73",
   375 => x"0b0b0b92",
   376 => x"882effaa",
   377 => x"388af004",
   378 => x"76880c02",
   379 => x"80c0050d",
   380 => x"0402f805",
   381 => x"0d7352c0",
   382 => x"0870882a",
   383 => x"70810651",
   384 => x"51517080",
   385 => x"2ef13871",
   386 => x"c00c7188",
   387 => x"0c028805",
   388 => x"0d0402e8",
   389 => x"050d8078",
   390 => x"57557570",
   391 => x"84055708",
   392 => x"53805472",
   393 => x"982a7388",
   394 => x"2b545271",
   395 => x"802ea238",
   396 => x"c0087088",
   397 => x"2a708106",
   398 => x"51515170",
   399 => x"802ef138",
   400 => x"71c00c81",
   401 => x"15811555",
   402 => x"55837425",
   403 => x"d63871ca",
   404 => x"3874880c",
   405 => x"0298050d",
   406 => x"0402ec05",
   407 => x"0d805184",
   408 => x"80800bfc",
   409 => x"800c8111",
   410 => x"70525584",
   411 => x"80805380",
   412 => x"5484fe52",
   413 => x"81117083",
   414 => x"ffff0670",
   415 => x"75708405",
   416 => x"570cfe14",
   417 => x"54515171",
   418 => x"8025e938",
   419 => x"81145483",
   420 => x"df7425dd",
   421 => x"38811551",
   422 => x"8ce60494",
   423 => x"0802940c",
   424 => x"fd3d0d80",
   425 => x"5394088c",
   426 => x"05085294",
   427 => x"08880508",
   428 => x"5182de3f",
   429 => x"88087088",
   430 => x"0c54853d",
   431 => x"0d940c04",
   432 => x"94080294",
   433 => x"0cfd3d0d",
   434 => x"81539408",
   435 => x"8c050852",
   436 => x"94088805",
   437 => x"085182b9",
   438 => x"3f880870",
   439 => x"880c5485",
   440 => x"3d0d940c",
   441 => x"04940802",
   442 => x"940cf93d",
   443 => x"0d800b94",
   444 => x"08fc050c",
   445 => x"94088805",
   446 => x"088025ab",
   447 => x"38940888",
   448 => x"05083094",
   449 => x"0888050c",
   450 => x"800b9408",
   451 => x"f4050c94",
   452 => x"08fc0508",
   453 => x"8838810b",
   454 => x"9408f405",
   455 => x"0c9408f4",
   456 => x"05089408",
   457 => x"fc050c94",
   458 => x"088c0508",
   459 => x"8025ab38",
   460 => x"94088c05",
   461 => x"08309408",
   462 => x"8c050c80",
   463 => x"0b9408f0",
   464 => x"050c9408",
   465 => x"fc050888",
   466 => x"38810b94",
   467 => x"08f0050c",
   468 => x"9408f005",
   469 => x"089408fc",
   470 => x"050c8053",
   471 => x"94088c05",
   472 => x"08529408",
   473 => x"88050851",
   474 => x"81a73f88",
   475 => x"08709408",
   476 => x"f8050c54",
   477 => x"9408fc05",
   478 => x"08802e8c",
   479 => x"389408f8",
   480 => x"05083094",
   481 => x"08f8050c",
   482 => x"9408f805",
   483 => x"0870880c",
   484 => x"54893d0d",
   485 => x"940c0494",
   486 => x"0802940c",
   487 => x"fb3d0d80",
   488 => x"0b9408fc",
   489 => x"050c9408",
   490 => x"88050880",
   491 => x"25933894",
   492 => x"08880508",
   493 => x"30940888",
   494 => x"050c810b",
   495 => x"9408fc05",
   496 => x"0c94088c",
   497 => x"05088025",
   498 => x"8c389408",
   499 => x"8c050830",
   500 => x"94088c05",
   501 => x"0c815394",
   502 => x"088c0508",
   503 => x"52940888",
   504 => x"050851ad",
   505 => x"3f880870",
   506 => x"9408f805",
   507 => x"0c549408",
   508 => x"fc050880",
   509 => x"2e8c3894",
   510 => x"08f80508",
   511 => x"309408f8",
   512 => x"050c9408",
   513 => x"f8050870",
   514 => x"880c5487",
   515 => x"3d0d940c",
   516 => x"04940802",
   517 => x"940cfd3d",
   518 => x"0d810b94",
   519 => x"08fc050c",
   520 => x"800b9408",
   521 => x"f8050c94",
   522 => x"088c0508",
   523 => x"94088805",
   524 => x"0827ac38",
   525 => x"9408fc05",
   526 => x"08802ea3",
   527 => x"38800b94",
   528 => x"088c0508",
   529 => x"24993894",
   530 => x"088c0508",
   531 => x"1094088c",
   532 => x"050c9408",
   533 => x"fc050810",
   534 => x"9408fc05",
   535 => x"0cc93994",
   536 => x"08fc0508",
   537 => x"802e80c9",
   538 => x"3894088c",
   539 => x"05089408",
   540 => x"88050826",
   541 => x"a1389408",
   542 => x"88050894",
   543 => x"088c0508",
   544 => x"31940888",
   545 => x"050c9408",
   546 => x"f8050894",
   547 => x"08fc0508",
   548 => x"079408f8",
   549 => x"050c9408",
   550 => x"fc050881",
   551 => x"2a9408fc",
   552 => x"050c9408",
   553 => x"8c050881",
   554 => x"2a94088c",
   555 => x"050cffaf",
   556 => x"39940890",
   557 => x"0508802e",
   558 => x"8f389408",
   559 => x"88050870",
   560 => x"9408f405",
   561 => x"0c518d39",
   562 => x"9408f805",
   563 => x"08709408",
   564 => x"f4050c51",
   565 => x"9408f405",
   566 => x"08880c85",
   567 => x"3d0d940c",
   568 => x"04000000",
   569 => x"00ffffff",
   570 => x"ff00ffff",
   571 => x"ffff00ff",
   572 => x"ffffff00",
   573 => x"30313233",
   574 => x"34353637",
   575 => x"38394142",
   576 => x"43444546",
   577 => x"00444546",
	others => x"00000000"
);

begin

process (clk)
begin
	if (clk'event and clk = '1') then
		if (from_zpu.memAWriteEnable = '1') and (from_zpu.memBWriteEnable = '1') and (from_zpu.memAAddr=from_zpu.memBAddr) and (from_zpu.memAWrite/=from_zpu.memBWrite) then
			report "write collision" severity failure;
		end if;
	
		if (from_zpu.memAWriteEnable = '1') then
			ram(to_integer(unsigned(from_zpu.memAAddr(maxAddrBitBRAM downto 2)))) := from_zpu.memAWrite;
			to_zpu.memARead <= from_zpu.memAWrite;
		else
			to_zpu.memARead <= ram(to_integer(unsigned(from_zpu.memAAddr(maxAddrBitBRAM downto 2))));
		end if;
	end if;
end process;

process (clk)
begin
	if (clk'event and clk = '1') then
		if (from_zpu.memBWriteEnable = '1') then
			ram(to_integer(unsigned(from_zpu.memBAddr(maxAddrBitBRAM downto 2)))) := from_zpu.memBWrite;
			to_zpu.memBRead <= from_zpu.memBWrite;
		else
			to_zpu.memBRead <= ram(to_integer(unsigned(from_zpu.memBAddr(maxAddrBitBRAM downto 2))));
		end if;
	end if;
end process;


end arch;

