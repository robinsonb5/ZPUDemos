-- ZPU
--
-- Copyright 2004-2008 oharboe - �yvind Harboe - oyvind.harboe@zylin.com
-- Modified by Alastair M. Robinson for the ZPUFlex project.
--
-- The FreeBSD license
-- 
-- Redistribution and use in source and binary forms, with or without
-- modification, are permitted provided that the following conditions
-- are met:
-- 
-- 1. Redistributions of source code must retain the above copyright
--    notice, this list of conditions and the following disclaimer.
-- 2. Redistributions in binary form must reproduce the above
--    copyright notice, this list of conditions and the following
--    disclaimer in the documentation and/or other materials
--    provided with the distribution.
-- 
-- THIS SOFTWARE IS PROVIDED BY THE ZPU PROJECT ``AS IS'' AND ANY
-- EXPRESS OR IMPLIED WARRANTIES, INCLUDING, BUT NOT LIMITED TO,
-- THE IMPLIED WARRANTIES OF MERCHANTABILITY AND FITNESS FOR A
-- PARTICULAR PURPOSE ARE DISCLAIMED. IN NO EVENT SHALL THE
-- ZPU PROJECT OR CONTRIBUTORS BE LIABLE FOR ANY DIRECT,
-- INDIRECT, INCIDENTAL, SPECIAL, EXEMPLARY, OR CONSEQUENTIAL DAMAGES
-- (INCLUDING, BUT NOT LIMITED TO, PROCUREMENT OF SUBSTITUTE GOODS
-- OR SERVICES; LOSS OF USE, DATA, OR PROFITS; OR BUSINESS INTERRUPTION)
-- HOWEVER CAUSED AND ON ANY THEORY OF LIABILITY, WHETHER IN CONTRACT,
-- STRICT LIABILITY, OR TORT (INCLUDING NEGLIGENCE OR OTHERWISE)
-- ARISING IN ANY WAY OUT OF THE USE OF THIS SOFTWARE, EVEN IF
-- ADVISED OF THE POSSIBILITY OF SUCH DAMAGE.
-- 
-- The views and conclusions contained in the software and documentation
-- are those of the authors and should not be interpreted as representing
-- official policies, either expressed or implied, of the ZPU Project.

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;


library work;
use work.zpupkg.all;

entity SDBootstrap_ROM is
generic
	(
		maxAddrBitBRAM : integer := maxAddrBitBRAMLimit -- Specify your actual ROM size to save LEs and unnecessary block RAM usage.
	);
port (
	clk : in std_logic;
	areset : in std_logic := '0';
	from_zpu : in ZPU_ToROM;
	to_zpu : out ZPU_FromROM
);
end SDBootstrap_ROM;

architecture arch of SDBootstrap_ROM is

type ram_type is array(natural range 0 to ((2**(maxAddrBitBRAM+1))/4)-1) of std_logic_vector(wordSize-1 downto 0);

shared variable ram : ram_type :=
(
     0 => x"84808080",
     1 => x"8c0b8480",
     2 => x"8081e004",
     3 => x"00848080",
     4 => x"808c04ff",
     5 => x"0d800404",
     6 => x"40000017",
     7 => x"00000000",
     8 => x"0b83ffe0",
     9 => x"80080b83",
    10 => x"ffe08408",
    11 => x"0b83ffe0",
    12 => x"88088480",
    13 => x"80809808",
    14 => x"2d0b83ff",
    15 => x"e0880c0b",
    16 => x"83ffe084",
    17 => x"0c0b83ff",
    18 => x"e0800c04",
    19 => x"00000000",
    20 => x"00000000",
    21 => x"00000000",
    22 => x"00000000",
    23 => x"00000000",
    24 => x"71fd0608",
    25 => x"72830609",
    26 => x"81058205",
    27 => x"832b2a83",
    28 => x"ffff0652",
    29 => x"0471fc06",
    30 => x"08728306",
    31 => x"09810583",
    32 => x"05101010",
    33 => x"2a81ff06",
    34 => x"520471fd",
    35 => x"060883ff",
    36 => x"ff738306",
    37 => x"09810582",
    38 => x"05832b2b",
    39 => x"09067383",
    40 => x"ffff0673",
    41 => x"83060981",
    42 => x"05820583",
    43 => x"2b0b2b07",
    44 => x"72fc060c",
    45 => x"51510471",
    46 => x"fc060884",
    47 => x"8080a5a0",
    48 => x"73830610",
    49 => x"10050806",
    50 => x"7381ff06",
    51 => x"73830609",
    52 => x"81058305",
    53 => x"1010102b",
    54 => x"0772fc06",
    55 => x"0c515104",
    56 => x"83ffe080",
    57 => x"7083fff6",
    58 => x"8c278e38",
    59 => x"80717084",
    60 => x"05530c84",
    61 => x"808081e4",
    62 => x"04848080",
    63 => x"808c5184",
    64 => x"80809388",
    65 => x"0402ec05",
    66 => x"0d765380",
    67 => x"5572752e",
    68 => x"be388754",
    69 => x"729c2a73",
    70 => x"842b5452",
    71 => x"71802e83",
    72 => x"38815589",
    73 => x"72258a38",
    74 => x"b7125284",
    75 => x"808082b4",
    76 => x"04b01252",
    77 => x"74802e89",
    78 => x"38715184",
    79 => x"808085a1",
    80 => x"2dff1454",
    81 => x"738025cc",
    82 => x"38848080",
    83 => x"82d704b0",
    84 => x"51848080",
    85 => x"85a12d80",
    86 => x"0b83ffe0",
    87 => x"800c0294",
    88 => x"050d0402",
    89 => x"c0050d02",
    90 => x"80c40557",
    91 => x"80707870",
    92 => x"84055a08",
    93 => x"72415f5d",
    94 => x"587c7084",
    95 => x"055e085a",
    96 => x"805b7998",
    97 => x"2a7a882b",
    98 => x"5b567589",
    99 => x"38775f84",
   100 => x"80808595",
   101 => x"047d802e",
   102 => x"81d33880",
   103 => x"5e7580e4",
   104 => x"2e8a3875",
   105 => x"80f82e09",
   106 => x"81068938",
   107 => x"76841871",
   108 => x"085e5854",
   109 => x"7580e42e",
   110 => x"a6387580",
   111 => x"e4268e38",
   112 => x"7580e32e",
   113 => x"80d93884",
   114 => x"808084ad",
   115 => x"047580f3",
   116 => x"2eb53875",
   117 => x"80f82e8f",
   118 => x"38848080",
   119 => x"84ad048a",
   120 => x"53848080",
   121 => x"83e90490",
   122 => x"5383ffe0",
   123 => x"e0527b51",
   124 => x"84808082",
   125 => x"852d83ff",
   126 => x"e0800883",
   127 => x"ffe0e05a",
   128 => x"55848080",
   129 => x"84c60476",
   130 => x"84187108",
   131 => x"70545b58",
   132 => x"54848080",
   133 => x"85c52d80",
   134 => x"55848080",
   135 => x"84c60476",
   136 => x"84187108",
   137 => x"58585484",
   138 => x"808084fd",
   139 => x"04a55184",
   140 => x"808085a1",
   141 => x"2d755184",
   142 => x"808085a1",
   143 => x"2d821858",
   144 => x"84808085",
   145 => x"880474ff",
   146 => x"16565480",
   147 => x"7425b938",
   148 => x"78708105",
   149 => x"5a848080",
   150 => x"80f52d70",
   151 => x"52568480",
   152 => x"8085a12d",
   153 => x"81185884",
   154 => x"808084c6",
   155 => x"0475a52e",
   156 => x"09810689",
   157 => x"38815e84",
   158 => x"80808588",
   159 => x"04755184",
   160 => x"808085a1",
   161 => x"2d811858",
   162 => x"811b5b83",
   163 => x"7b25fdf2",
   164 => x"3875fde5",
   165 => x"387e83ff",
   166 => x"e0800c02",
   167 => x"80c0050d",
   168 => x"0402f805",
   169 => x"0d7352c0",
   170 => x"0870882a",
   171 => x"70810651",
   172 => x"51517080",
   173 => x"2ef13871",
   174 => x"c00c7183",
   175 => x"ffe0800c",
   176 => x"0288050d",
   177 => x"0402e805",
   178 => x"0d807857",
   179 => x"55757084",
   180 => x"05570853",
   181 => x"80547298",
   182 => x"2a73882b",
   183 => x"54527180",
   184 => x"2ea238c0",
   185 => x"0870882a",
   186 => x"70810651",
   187 => x"51517080",
   188 => x"2ef13871",
   189 => x"c00c8115",
   190 => x"81155555",
   191 => x"837425d6",
   192 => x"3871ca38",
   193 => x"7483ffe0",
   194 => x"800c0298",
   195 => x"050d0402",
   196 => x"f4050dd4",
   197 => x"5281ff72",
   198 => x"0c710853",
   199 => x"81ff720c",
   200 => x"72882b83",
   201 => x"fe800672",
   202 => x"087081ff",
   203 => x"06515253",
   204 => x"81ff720c",
   205 => x"72710788",
   206 => x"2b720870",
   207 => x"81ff0651",
   208 => x"525381ff",
   209 => x"720c7271",
   210 => x"07882b72",
   211 => x"087081ff",
   212 => x"06720783",
   213 => x"ffe0800c",
   214 => x"5253028c",
   215 => x"050d0402",
   216 => x"f4050d74",
   217 => x"767181ff",
   218 => x"06d40c53",
   219 => x"5383fff1",
   220 => x"a0088538",
   221 => x"71892b52",
   222 => x"71982ad4",
   223 => x"0c71902a",
   224 => x"7081ff06",
   225 => x"d40c5171",
   226 => x"882a7081",
   227 => x"ff06d40c",
   228 => x"517181ff",
   229 => x"06d40c72",
   230 => x"902a7081",
   231 => x"ff06d40c",
   232 => x"51d40870",
   233 => x"81ff0651",
   234 => x"5182b8bf",
   235 => x"527081ff",
   236 => x"2e098106",
   237 => x"943881ff",
   238 => x"0bd40cd4",
   239 => x"087081ff",
   240 => x"06ff1454",
   241 => x"515171e5",
   242 => x"387083ff",
   243 => x"e0800c02",
   244 => x"8c050d04",
   245 => x"02fc050d",
   246 => x"81c75181",
   247 => x"ff0bd40c",
   248 => x"ff115170",
   249 => x"8025f438",
   250 => x"0284050d",
   251 => x"0402f005",
   252 => x"0d848080",
   253 => x"87d42d81",
   254 => x"9c9f5380",
   255 => x"5287fc80",
   256 => x"f7518480",
   257 => x"8086df2d",
   258 => x"83ffe080",
   259 => x"085483ff",
   260 => x"e0800881",
   261 => x"2e098106",
   262 => x"ae3881ff",
   263 => x"0bd40c82",
   264 => x"0a52849c",
   265 => x"80e95184",
   266 => x"808086df",
   267 => x"2d83ffe0",
   268 => x"80088e38",
   269 => x"81ff0bd4",
   270 => x"0c735384",
   271 => x"808088ce",
   272 => x"04848080",
   273 => x"87d42dff",
   274 => x"135372ff",
   275 => x"ae387283",
   276 => x"ffe0800c",
   277 => x"0290050d",
   278 => x"0402f405",
   279 => x"0d81ff0b",
   280 => x"d40c8480",
   281 => x"80a5b051",
   282 => x"84808085",
   283 => x"c52d9353",
   284 => x"805287fc",
   285 => x"80c15184",
   286 => x"808086df",
   287 => x"2d83ffe0",
   288 => x"80088e38",
   289 => x"81ff0bd4",
   290 => x"0c815384",
   291 => x"8080899d",
   292 => x"04848080",
   293 => x"87d42dff",
   294 => x"135372d4",
   295 => x"387283ff",
   296 => x"e0800c02",
   297 => x"8c050d04",
   298 => x"02f0050d",
   299 => x"84808087",
   300 => x"d42d83aa",
   301 => x"52849c80",
   302 => x"c8518480",
   303 => x"8086df2d",
   304 => x"83ffe080",
   305 => x"0883ffe0",
   306 => x"80085384",
   307 => x"8080a5bc",
   308 => x"52538480",
   309 => x"8082e32d",
   310 => x"72812e09",
   311 => x"8106a938",
   312 => x"84808086",
   313 => x"8f2d83ff",
   314 => x"e0800883",
   315 => x"ffff0653",
   316 => x"7283aa2e",
   317 => x"bb3883ff",
   318 => x"e0800852",
   319 => x"848080a5",
   320 => x"d4518480",
   321 => x"8082e32d",
   322 => x"84808088",
   323 => x"d92d8480",
   324 => x"808aa804",
   325 => x"81548480",
   326 => x"808bd304",
   327 => x"848080a5",
   328 => x"ec518480",
   329 => x"8082e32d",
   330 => x"80548480",
   331 => x"808bd304",
   332 => x"81ff0bd4",
   333 => x"0cb15384",
   334 => x"808087ed",
   335 => x"2d83ffe0",
   336 => x"8008802e",
   337 => x"80fe3880",
   338 => x"5287fc80",
   339 => x"fa518480",
   340 => x"8086df2d",
   341 => x"83ffe080",
   342 => x"0880d738",
   343 => x"83ffe080",
   344 => x"08528480",
   345 => x"80a68851",
   346 => x"84808082",
   347 => x"e32d81ff",
   348 => x"0bd40cd4",
   349 => x"087081ff",
   350 => x"06705484",
   351 => x"8080a694",
   352 => x"53515384",
   353 => x"808082e3",
   354 => x"2d81ff0b",
   355 => x"d40c81ff",
   356 => x"0bd40c81",
   357 => x"ff0bd40c",
   358 => x"81ff0bd4",
   359 => x"0c72862a",
   360 => x"70810670",
   361 => x"56515372",
   362 => x"802ea838",
   363 => x"8480808a",
   364 => x"940483ff",
   365 => x"e0800852",
   366 => x"848080a6",
   367 => x"88518480",
   368 => x"8082e32d",
   369 => x"72822efe",
   370 => x"d338ff13",
   371 => x"5372fee7",
   372 => x"38725473",
   373 => x"83ffe080",
   374 => x"0c029005",
   375 => x"0d0402f4",
   376 => x"050d810b",
   377 => x"83fff1a0",
   378 => x"0cd00870",
   379 => x"8f2a7081",
   380 => x"06515153",
   381 => x"72f33872",
   382 => x"d00c8480",
   383 => x"8087d42d",
   384 => x"848080a6",
   385 => x"a4518480",
   386 => x"8085c52d",
   387 => x"d008708f",
   388 => x"2a708106",
   389 => x"51515372",
   390 => x"f338810b",
   391 => x"d00c8753",
   392 => x"805284d4",
   393 => x"80c05184",
   394 => x"808086df",
   395 => x"2d83ffe0",
   396 => x"8008812e",
   397 => x"97387282",
   398 => x"2e098106",
   399 => x"89388053",
   400 => x"8480808d",
   401 => x"8d04ff13",
   402 => x"5372d538",
   403 => x"84808089",
   404 => x"a82d83ff",
   405 => x"e0800883",
   406 => x"fff1a00c",
   407 => x"83ffe080",
   408 => x"088e3881",
   409 => x"5287fc80",
   410 => x"d0518480",
   411 => x"8086df2d",
   412 => x"81ff0bd4",
   413 => x"0cd00870",
   414 => x"8f2a7081",
   415 => x"06515153",
   416 => x"72f33872",
   417 => x"d00c81ff",
   418 => x"0bd40c81",
   419 => x"537283ff",
   420 => x"e0800c02",
   421 => x"8c050d04",
   422 => x"800b83ff",
   423 => x"e0800c04",
   424 => x"02e0050d",
   425 => x"797b5757",
   426 => x"805881ff",
   427 => x"0bd40cd0",
   428 => x"08708f2a",
   429 => x"70810651",
   430 => x"515473f3",
   431 => x"3882810b",
   432 => x"d00c81ff",
   433 => x"0bd40c76",
   434 => x"5287fc80",
   435 => x"d1518480",
   436 => x"8086df2d",
   437 => x"80dbc6df",
   438 => x"5583ffe0",
   439 => x"8008802e",
   440 => x"9b3883ff",
   441 => x"e0800853",
   442 => x"76528480",
   443 => x"80a6b051",
   444 => x"84808082",
   445 => x"e32d8480",
   446 => x"808ed204",
   447 => x"81ff0bd4",
   448 => x"0cd40870",
   449 => x"81ff0651",
   450 => x"547381fe",
   451 => x"2e098106",
   452 => x"a53880ff",
   453 => x"54848080",
   454 => x"868f2d83",
   455 => x"ffe08008",
   456 => x"76708405",
   457 => x"580cff14",
   458 => x"54738025",
   459 => x"e8388158",
   460 => x"8480808e",
   461 => x"bc04ff15",
   462 => x"5574c138",
   463 => x"81ff0bd4",
   464 => x"0cd00870",
   465 => x"8f2a7081",
   466 => x"06515154",
   467 => x"73f33873",
   468 => x"d00c7783",
   469 => x"ffe0800c",
   470 => x"02a0050d",
   471 => x"0402f405",
   472 => x"0d747088",
   473 => x"2a83fe80",
   474 => x"06707298",
   475 => x"2a077288",
   476 => x"2b87fc80",
   477 => x"80067398",
   478 => x"2b81f00a",
   479 => x"06717307",
   480 => x"0783ffe0",
   481 => x"800c5651",
   482 => x"5351028c",
   483 => x"050d0402",
   484 => x"f8050d02",
   485 => x"8e058480",
   486 => x"8080f52d",
   487 => x"74882b07",
   488 => x"7083ffff",
   489 => x"0683ffe0",
   490 => x"800c5102",
   491 => x"88050d04",
   492 => x"02f8050d",
   493 => x"7370902b",
   494 => x"71902a07",
   495 => x"83ffe080",
   496 => x"0c520288",
   497 => x"050d0402",
   498 => x"fc050d73",
   499 => x"81df06c9",
   500 => x"05517080",
   501 => x"258438a7",
   502 => x"11517284",
   503 => x"2b710783",
   504 => x"ffe0800c",
   505 => x"0284050d",
   506 => x"0402f005",
   507 => x"0d029705",
   508 => x"84808080",
   509 => x"f52d83ff",
   510 => x"f1c00881",
   511 => x"0583fff1",
   512 => x"c00c5473",
   513 => x"80d32e09",
   514 => x"8106a338",
   515 => x"800b83ff",
   516 => x"f1c00c80",
   517 => x"0b83fff1",
   518 => x"b00c800b",
   519 => x"83fff1c4",
   520 => x"0c800b83",
   521 => x"fff1ac0c",
   522 => x"84808093",
   523 => x"830483ff",
   524 => x"f1c00852",
   525 => x"71812e09",
   526 => x"8106bc38",
   527 => x"83fff1ac",
   528 => x"087481df",
   529 => x"06c90552",
   530 => x"52708025",
   531 => x"8438a711",
   532 => x"5171842b",
   533 => x"71077083",
   534 => x"fff1ac0c",
   535 => x"70525283",
   536 => x"72258538",
   537 => x"8a723151",
   538 => x"70108205",
   539 => x"83fff1b8",
   540 => x"0c848080",
   541 => x"93830471",
   542 => x"8324a638",
   543 => x"83fff1c4",
   544 => x"087481df",
   545 => x"06c90552",
   546 => x"52708025",
   547 => x"8438a711",
   548 => x"5171842b",
   549 => x"710783ff",
   550 => x"f1c40c84",
   551 => x"80809383",
   552 => x"0483fff1",
   553 => x"b8088305",
   554 => x"51717124",
   555 => x"a63883ff",
   556 => x"f1b00874",
   557 => x"81df06c9",
   558 => x"05525270",
   559 => x"80258438",
   560 => x"a7115171",
   561 => x"842b7107",
   562 => x"83fff1b0",
   563 => x"0c848080",
   564 => x"92c20483",
   565 => x"fff1ac08",
   566 => x"ff115253",
   567 => x"70822681",
   568 => x"973883ff",
   569 => x"f1c40810",
   570 => x"81055171",
   571 => x"712480df",
   572 => x"3883fff1",
   573 => x"bc087481",
   574 => x"df06c905",
   575 => x"52527080",
   576 => x"258438a7",
   577 => x"11517184",
   578 => x"2b710770",
   579 => x"83fff1bc",
   580 => x"0c83fff1",
   581 => x"b408ff05",
   582 => x"83fff1b4",
   583 => x"0c5283ff",
   584 => x"f1b40880",
   585 => x"2580dc38",
   586 => x"83fff1b0",
   587 => x"08517171",
   588 => x"84808081",
   589 => x"b72d83ff",
   590 => x"f1b00881",
   591 => x"0583fff1",
   592 => x"b00c810b",
   593 => x"83fff1b4",
   594 => x"0c848080",
   595 => x"93830483",
   596 => x"fff1b408",
   597 => x"ae3883ff",
   598 => x"f1bc0884",
   599 => x"2b7083ff",
   600 => x"f1bc0c83",
   601 => x"fff1b008",
   602 => x"52527171",
   603 => x"84808081",
   604 => x"b72d8480",
   605 => x"80938304",
   606 => x"86732587",
   607 => x"38848080",
   608 => x"80932d02",
   609 => x"90050d04",
   610 => x"02ec050d",
   611 => x"800bfc80",
   612 => x"0c848080",
   613 => x"a6d05184",
   614 => x"808085c5",
   615 => x"2d848080",
   616 => x"8bde2d83",
   617 => x"ffe08008",
   618 => x"802e8286",
   619 => x"38848080",
   620 => x"a6e85184",
   621 => x"808085c5",
   622 => x"2d848080",
   623 => x"96c82d83",
   624 => x"ffe1a052",
   625 => x"848080a7",
   626 => x"80518480",
   627 => x"80a3fe2d",
   628 => x"83ffe080",
   629 => x"08802e81",
   630 => x"cd3883ff",
   631 => x"e1a00b84",
   632 => x"8080a78c",
   633 => x"52548480",
   634 => x"8085c52d",
   635 => x"80557370",
   636 => x"81055584",
   637 => x"808080f5",
   638 => x"2d5372a0",
   639 => x"2e80e638",
   640 => x"72c00c72",
   641 => x"a32e8184",
   642 => x"387280c7",
   643 => x"2e098106",
   644 => x"8d388480",
   645 => x"8080932d",
   646 => x"84808094",
   647 => x"c004728a",
   648 => x"2e098106",
   649 => x"8d388480",
   650 => x"80808c2d",
   651 => x"84808094",
   652 => x"c0047280",
   653 => x"cc2e0981",
   654 => x"06863883",
   655 => x"ffe1a054",
   656 => x"7281df06",
   657 => x"f0057081",
   658 => x"ff065153",
   659 => x"b8732789",
   660 => x"38ef1370",
   661 => x"81ff0651",
   662 => x"5374842b",
   663 => x"73075584",
   664 => x"808093ee",
   665 => x"0472a32e",
   666 => x"a3387370",
   667 => x"81055584",
   668 => x"808080f5",
   669 => x"2d5372a0",
   670 => x"2ef038ff",
   671 => x"14755370",
   672 => x"52548480",
   673 => x"80a3fe2d",
   674 => x"74fc800c",
   675 => x"73708105",
   676 => x"55848080",
   677 => x"80f52d53",
   678 => x"728a2e09",
   679 => x"8106ed38",
   680 => x"84808093",
   681 => x"ec048480",
   682 => x"80a7a051",
   683 => x"84808085",
   684 => x"c52d8480",
   685 => x"80a7bc51",
   686 => x"84808085",
   687 => x"c52dae51",
   688 => x"84808085",
   689 => x"a12dbd84",
   690 => x"bf55c008",
   691 => x"70892a70",
   692 => x"81065154",
   693 => x"5472802e",
   694 => x"92387381",
   695 => x"ff065184",
   696 => x"80808fe9",
   697 => x"2d848080",
   698 => x"95c604ff",
   699 => x"155574ff",
   700 => x"2e098106",
   701 => x"d5388480",
   702 => x"8095be04",
   703 => x"02e8050d",
   704 => x"77797b58",
   705 => x"55558053",
   706 => x"727625af",
   707 => x"38747081",
   708 => x"05568480",
   709 => x"8080f52d",
   710 => x"74708105",
   711 => x"56848080",
   712 => x"80f52d52",
   713 => x"5271712e",
   714 => x"89388151",
   715 => x"84808096",
   716 => x"bd048113",
   717 => x"53848080",
   718 => x"96880480",
   719 => x"517083ff",
   720 => x"e0800c02",
   721 => x"98050d04",
   722 => x"02d8050d",
   723 => x"800b83ff",
   724 => x"f5f80c84",
   725 => x"8080a7d0",
   726 => x"51848080",
   727 => x"85c52d83",
   728 => x"fff1d452",
   729 => x"80518480",
   730 => x"808da02d",
   731 => x"83ffe080",
   732 => x"085483ff",
   733 => x"e0800895",
   734 => x"38848080",
   735 => x"a7e05184",
   736 => x"808085c5",
   737 => x"2d735584",
   738 => x"80809ef7",
   739 => x"04848080",
   740 => x"a7f45184",
   741 => x"808085c5",
   742 => x"2d805681",
   743 => x"0b83fff1",
   744 => x"c80c8853",
   745 => x"848080a8",
   746 => x"8c5283ff",
   747 => x"f28a5184",
   748 => x"808095fc",
   749 => x"2d83ffe0",
   750 => x"8008762e",
   751 => x"0981068b",
   752 => x"3883ffe0",
   753 => x"800883ff",
   754 => x"f1c80c88",
   755 => x"53848080",
   756 => x"a8985283",
   757 => x"fff2a651",
   758 => x"84808095",
   759 => x"fc2d83ff",
   760 => x"e080088b",
   761 => x"3883ffe0",
   762 => x"800883ff",
   763 => x"f1c80c83",
   764 => x"fff1c808",
   765 => x"52848080",
   766 => x"a8a45184",
   767 => x"808082e3",
   768 => x"2d83fff1",
   769 => x"c808802e",
   770 => x"81cb3883",
   771 => x"fff59a0b",
   772 => x"84808080",
   773 => x"f52d83ff",
   774 => x"f59b0b84",
   775 => x"808080f5",
   776 => x"2d71982b",
   777 => x"71902b07",
   778 => x"83fff59c",
   779 => x"0b848080",
   780 => x"80f52d70",
   781 => x"882b7207",
   782 => x"83fff59d",
   783 => x"0b848080",
   784 => x"80f52d71",
   785 => x"0783fff5",
   786 => x"d20b8480",
   787 => x"8080f52d",
   788 => x"83fff5d3",
   789 => x"0b848080",
   790 => x"80f52d71",
   791 => x"882b0753",
   792 => x"5f54525a",
   793 => x"56575573",
   794 => x"81abaa2e",
   795 => x"09810695",
   796 => x"38755184",
   797 => x"80808edd",
   798 => x"2d83ffe0",
   799 => x"80085684",
   800 => x"8080999e",
   801 => x"047382d4",
   802 => x"d52e9338",
   803 => x"848080a8",
   804 => x"b8518480",
   805 => x"8085c52d",
   806 => x"8480809b",
   807 => x"aa047552",
   808 => x"848080a8",
   809 => x"d8518480",
   810 => x"8082e32d",
   811 => x"83fff1d4",
   812 => x"52755184",
   813 => x"80808da0",
   814 => x"2d83ffe0",
   815 => x"80085583",
   816 => x"ffe08008",
   817 => x"802e85af",
   818 => x"38848080",
   819 => x"a8f05184",
   820 => x"808085c5",
   821 => x"2d848080",
   822 => x"a9985184",
   823 => x"808082e3",
   824 => x"2d885384",
   825 => x"8080a898",
   826 => x"5283fff2",
   827 => x"a6518480",
   828 => x"8095fc2d",
   829 => x"83ffe080",
   830 => x"088e3881",
   831 => x"0b83fff5",
   832 => x"f80c8480",
   833 => x"809ab604",
   834 => x"88538480",
   835 => x"80a88c52",
   836 => x"83fff28a",
   837 => x"51848080",
   838 => x"95fc2d83",
   839 => x"ffe08008",
   840 => x"802e9338",
   841 => x"848080a9",
   842 => x"b0518480",
   843 => x"8082e32d",
   844 => x"8480809b",
   845 => x"aa0483ff",
   846 => x"f5d20b84",
   847 => x"808080f5",
   848 => x"2d547380",
   849 => x"d52e0981",
   850 => x"0680df38",
   851 => x"83fff5d3",
   852 => x"0b848080",
   853 => x"80f52d54",
   854 => x"7381aa2e",
   855 => x"09810680",
   856 => x"c938800b",
   857 => x"83fff1d4",
   858 => x"0b848080",
   859 => x"80f52d56",
   860 => x"547481e9",
   861 => x"2e833881",
   862 => x"547481eb",
   863 => x"2e8c3880",
   864 => x"5573752e",
   865 => x"09810683",
   866 => x"ee3883ff",
   867 => x"f1df0b84",
   868 => x"808080f5",
   869 => x"2d597892",
   870 => x"3883fff1",
   871 => x"e00b8480",
   872 => x"8080f52d",
   873 => x"5473822e",
   874 => x"89388055",
   875 => x"8480809e",
   876 => x"f70483ff",
   877 => x"f1e10b84",
   878 => x"808080f5",
   879 => x"2d7083ff",
   880 => x"f6800cff",
   881 => x"117083ff",
   882 => x"f5f40c54",
   883 => x"52848080",
   884 => x"a9d05184",
   885 => x"808082e3",
   886 => x"2d83fff1",
   887 => x"e20b8480",
   888 => x"8080f52d",
   889 => x"83fff1e3",
   890 => x"0b848080",
   891 => x"80f52d56",
   892 => x"76057582",
   893 => x"80290570",
   894 => x"83fff5e8",
   895 => x"0c83fff1",
   896 => x"e40b8480",
   897 => x"8080f52d",
   898 => x"7083fff5",
   899 => x"e40c83ff",
   900 => x"f5f80859",
   901 => x"57587680",
   902 => x"2e81ec38",
   903 => x"88538480",
   904 => x"80a89852",
   905 => x"83fff2a6",
   906 => x"51848080",
   907 => x"95fc2d78",
   908 => x"5583ffe0",
   909 => x"800882bf",
   910 => x"3883fff6",
   911 => x"80087084",
   912 => x"2b83fff5",
   913 => x"d40c7083",
   914 => x"fff5fc0c",
   915 => x"83fff1f9",
   916 => x"0b848080",
   917 => x"80f52d83",
   918 => x"fff1f80b",
   919 => x"84808080",
   920 => x"f52d7182",
   921 => x"80290583",
   922 => x"fff1fa0b",
   923 => x"84808080",
   924 => x"f52d7084",
   925 => x"80802912",
   926 => x"83fff1fb",
   927 => x"0b848080",
   928 => x"80f52d70",
   929 => x"81800a29",
   930 => x"127083ff",
   931 => x"f1cc0c83",
   932 => x"fff5e408",
   933 => x"712983ff",
   934 => x"f5e80805",
   935 => x"7083fff6",
   936 => x"880c83ff",
   937 => x"f2810b84",
   938 => x"808080f5",
   939 => x"2d83fff2",
   940 => x"800b8480",
   941 => x"8080f52d",
   942 => x"71828029",
   943 => x"0583fff2",
   944 => x"820b8480",
   945 => x"8080f52d",
   946 => x"70848080",
   947 => x"291283ff",
   948 => x"f2830b84",
   949 => x"808080f5",
   950 => x"2d70982b",
   951 => x"81f00a06",
   952 => x"72057083",
   953 => x"fff1d00c",
   954 => x"fe117e29",
   955 => x"770583ff",
   956 => x"f5f00c52",
   957 => x"5752575d",
   958 => x"5751525f",
   959 => x"525c5757",
   960 => x"57848080",
   961 => x"9ef50483",
   962 => x"fff1e60b",
   963 => x"84808080",
   964 => x"f52d83ff",
   965 => x"f1e50b84",
   966 => x"808080f5",
   967 => x"2d718280",
   968 => x"29057083",
   969 => x"fff5d40c",
   970 => x"70a02983",
   971 => x"ff057089",
   972 => x"2a7083ff",
   973 => x"f5fc0c83",
   974 => x"fff1eb0b",
   975 => x"84808080",
   976 => x"f52d83ff",
   977 => x"f1ea0b84",
   978 => x"808080f5",
   979 => x"2d718280",
   980 => x"29057083",
   981 => x"fff1cc0c",
   982 => x"7b71291e",
   983 => x"7083fff5",
   984 => x"f00c7d83",
   985 => x"fff1d00c",
   986 => x"730583ff",
   987 => x"f6880c55",
   988 => x"5e515155",
   989 => x"55815574",
   990 => x"83ffe080",
   991 => x"0c02a805",
   992 => x"0d0402ec",
   993 => x"050d7670",
   994 => x"872c7180",
   995 => x"ff065556",
   996 => x"5483fff5",
   997 => x"f8088a38",
   998 => x"73882c74",
   999 => x"81ff0654",
  1000 => x"5583fff1",
  1001 => x"d45283ff",
  1002 => x"f5e80815",
  1003 => x"51848080",
  1004 => x"8da02d83",
  1005 => x"ffe08008",
  1006 => x"5483ffe0",
  1007 => x"8008802e",
  1008 => x"80c93883",
  1009 => x"fff5f808",
  1010 => x"802ea238",
  1011 => x"72842983",
  1012 => x"fff1d405",
  1013 => x"70085253",
  1014 => x"8480808e",
  1015 => x"dd2d83ff",
  1016 => x"e08008f0",
  1017 => x"0a065384",
  1018 => x"8080a089",
  1019 => x"04721083",
  1020 => x"fff1d405",
  1021 => x"70848080",
  1022 => x"80e02d52",
  1023 => x"53848080",
  1024 => x"8f8f2d83",
  1025 => x"ffe08008",
  1026 => x"53725473",
  1027 => x"83ffe080",
  1028 => x"0c029405",
  1029 => x"0d0402c8",
  1030 => x"050d7f61",
  1031 => x"5f5b800b",
  1032 => x"83fff1d0",
  1033 => x"0883fff5",
  1034 => x"f008595d",
  1035 => x"5683fff5",
  1036 => x"f808762e",
  1037 => x"8f3883ff",
  1038 => x"f6800884",
  1039 => x"2b588480",
  1040 => x"80a0cc04",
  1041 => x"83fff5fc",
  1042 => x"08842b58",
  1043 => x"80597878",
  1044 => x"2781dc38",
  1045 => x"788f06a0",
  1046 => x"17575473",
  1047 => x"963883ff",
  1048 => x"f1d45276",
  1049 => x"51811757",
  1050 => x"8480808d",
  1051 => x"a02d83ff",
  1052 => x"f1d45680",
  1053 => x"76848080",
  1054 => x"80f52d56",
  1055 => x"5474742e",
  1056 => x"83388154",
  1057 => x"7481e52e",
  1058 => x"819c3881",
  1059 => x"70750655",
  1060 => x"5d73802e",
  1061 => x"8190388b",
  1062 => x"16848080",
  1063 => x"80f52d98",
  1064 => x"065a7981",
  1065 => x"81388b53",
  1066 => x"7d527551",
  1067 => x"84808095",
  1068 => x"fc2d83ff",
  1069 => x"e0800880",
  1070 => x"ed389c16",
  1071 => x"08518480",
  1072 => x"808edd2d",
  1073 => x"83ffe080",
  1074 => x"08841c0c",
  1075 => x"9a168480",
  1076 => x"8080e02d",
  1077 => x"51848080",
  1078 => x"8f8f2d83",
  1079 => x"ffe08008",
  1080 => x"83ffe080",
  1081 => x"08881d0c",
  1082 => x"83ffe080",
  1083 => x"08555583",
  1084 => x"fff5f808",
  1085 => x"802ea038",
  1086 => x"94168480",
  1087 => x"8080e02d",
  1088 => x"51848080",
  1089 => x"8f8f2d83",
  1090 => x"ffe08008",
  1091 => x"902b83ff",
  1092 => x"f00a0670",
  1093 => x"16515473",
  1094 => x"881c0c79",
  1095 => x"7b0c7c54",
  1096 => x"848080a2",
  1097 => x"f7048119",
  1098 => x"59848080",
  1099 => x"a0ce0483",
  1100 => x"fff5f808",
  1101 => x"802ebe38",
  1102 => x"7b518480",
  1103 => x"809f822d",
  1104 => x"83ffe080",
  1105 => x"0883ffe0",
  1106 => x"800880ff",
  1107 => x"fffff806",
  1108 => x"555c7380",
  1109 => x"fffffff8",
  1110 => x"2e9b3883",
  1111 => x"ffe08008",
  1112 => x"fe0583ff",
  1113 => x"f6800829",
  1114 => x"83fff688",
  1115 => x"08055784",
  1116 => x"8080a0cc",
  1117 => x"04805473",
  1118 => x"83ffe080",
  1119 => x"0c02b805",
  1120 => x"0d0402f4",
  1121 => x"050d7470",
  1122 => x"08810571",
  1123 => x"0c700883",
  1124 => x"fff5f408",
  1125 => x"06535371",
  1126 => x"93388813",
  1127 => x"08518480",
  1128 => x"809f822d",
  1129 => x"83ffe080",
  1130 => x"0888140c",
  1131 => x"810b83ff",
  1132 => x"e0800c02",
  1133 => x"8c050d04",
  1134 => x"02f0050d",
  1135 => x"75881108",
  1136 => x"fe0583ff",
  1137 => x"f6800829",
  1138 => x"83fff688",
  1139 => x"08117208",
  1140 => x"83fff5f4",
  1141 => x"08060579",
  1142 => x"55535454",
  1143 => x"8480808d",
  1144 => x"a02d83ff",
  1145 => x"e0800853",
  1146 => x"83ffe080",
  1147 => x"08802e83",
  1148 => x"38815372",
  1149 => x"83ffe080",
  1150 => x"0c029005",
  1151 => x"0d0402ec",
  1152 => x"050d7678",
  1153 => x"715483ff",
  1154 => x"f5d85354",
  1155 => x"55848080",
  1156 => x"a0962d83",
  1157 => x"ffe08008",
  1158 => x"5483ffe0",
  1159 => x"8008802e",
  1160 => x"80ce3884",
  1161 => x"8080a9f4",
  1162 => x"51848080",
  1163 => x"85c52d83",
  1164 => x"fff5dc08",
  1165 => x"83ff0589",
  1166 => x"2a558054",
  1167 => x"73752580",
  1168 => x"d1387252",
  1169 => x"83fff5d8",
  1170 => x"51848080",
  1171 => x"a3b82d83",
  1172 => x"ffe08008",
  1173 => x"802eaf38",
  1174 => x"83fff5d8",
  1175 => x"51848080",
  1176 => x"a3822d84",
  1177 => x"80138115",
  1178 => x"55538480",
  1179 => x"80a4bc04",
  1180 => x"74528480",
  1181 => x"80aa9051",
  1182 => x"84808082",
  1183 => x"e32d7353",
  1184 => x"848080a5",
  1185 => x"940483ff",
  1186 => x"e0800853",
  1187 => x"848080a5",
  1188 => x"94048153",
  1189 => x"7283ffe0",
  1190 => x"800c0294",
  1191 => x"050d0400",
  1192 => x"00ffffff",
  1193 => x"ff00ffff",
  1194 => x"ffff00ff",
  1195 => x"ffffff00",
  1196 => x"436d645f",
  1197 => x"696e6974",
  1198 => x"0a000000",
  1199 => x"636d645f",
  1200 => x"434d4438",
  1201 => x"20726573",
  1202 => x"706f6e73",
  1203 => x"653a2025",
  1204 => x"640a0000",
  1205 => x"434d4438",
  1206 => x"5f342072",
  1207 => x"6573706f",
  1208 => x"6e73653a",
  1209 => x"2025640a",
  1210 => x"00000000",
  1211 => x"53444843",
  1212 => x"20496e69",
  1213 => x"7469616c",
  1214 => x"697a6174",
  1215 => x"696f6e20",
  1216 => x"6572726f",
  1217 => x"72210a00",
  1218 => x"434d4435",
  1219 => x"38202564",
  1220 => x"0a202000",
  1221 => x"434d4435",
  1222 => x"385f3220",
  1223 => x"25640a20",
  1224 => x"20000000",
  1225 => x"53504920",
  1226 => x"496e6974",
  1227 => x"28290a00",
  1228 => x"52656164",
  1229 => x"20636f6d",
  1230 => x"6d616e64",
  1231 => x"20666169",
  1232 => x"6c656420",
  1233 => x"61742025",
  1234 => x"64202825",
  1235 => x"64290a00",
  1236 => x"496e6974",
  1237 => x"69616c69",
  1238 => x"7a696e67",
  1239 => x"20534420",
  1240 => x"63617264",
  1241 => x"0a000000",
  1242 => x"48756e74",
  1243 => x"696e6720",
  1244 => x"666f7220",
  1245 => x"70617274",
  1246 => x"6974696f",
  1247 => x"6e0a0000",
  1248 => x"4d414e49",
  1249 => x"46455354",
  1250 => x"4d535400",
  1251 => x"50617273",
  1252 => x"696e6720",
  1253 => x"6d616e69",
  1254 => x"66657374",
  1255 => x"0a000000",
  1256 => x"4c6f6164",
  1257 => x"696e6720",
  1258 => x"6d616e69",
  1259 => x"66657374",
  1260 => x"20666169",
  1261 => x"6c65640a",
  1262 => x"00000000",
  1263 => x"426f6f74",
  1264 => x"696e6720",
  1265 => x"66726f6d",
  1266 => x"20525332",
  1267 => x"33322e00",
  1268 => x"52656164",
  1269 => x"696e6720",
  1270 => x"4d42520a",
  1271 => x"00000000",
  1272 => x"52656164",
  1273 => x"206f6620",
  1274 => x"4d425220",
  1275 => x"6661696c",
  1276 => x"65640a00",
  1277 => x"4d425220",
  1278 => x"73756363",
  1279 => x"65737366",
  1280 => x"756c6c79",
  1281 => x"20726561",
  1282 => x"640a0000",
  1283 => x"46415431",
  1284 => x"36202020",
  1285 => x"00000000",
  1286 => x"46415433",
  1287 => x"32202020",
  1288 => x"00000000",
  1289 => x"50617274",
  1290 => x"6974696f",
  1291 => x"6e636f75",
  1292 => x"6e742025",
  1293 => x"640a0000",
  1294 => x"4e6f2070",
  1295 => x"61727469",
  1296 => x"74696f6e",
  1297 => x"20736967",
  1298 => x"6e617475",
  1299 => x"72652066",
  1300 => x"6f756e64",
  1301 => x"0a000000",
  1302 => x"52656164",
  1303 => x"696e6720",
  1304 => x"626f6f74",
  1305 => x"20736563",
  1306 => x"746f7220",
  1307 => x"25640a00",
  1308 => x"52656164",
  1309 => x"20626f6f",
  1310 => x"74207365",
  1311 => x"63746f72",
  1312 => x"2066726f",
  1313 => x"6d206669",
  1314 => x"72737420",
  1315 => x"70617274",
  1316 => x"6974696f",
  1317 => x"6e0a0000",
  1318 => x"48756e74",
  1319 => x"696e6720",
  1320 => x"666f7220",
  1321 => x"66696c65",
  1322 => x"73797374",
  1323 => x"656d0a00",
  1324 => x"556e7375",
  1325 => x"70706f72",
  1326 => x"74656420",
  1327 => x"70617274",
  1328 => x"6974696f",
  1329 => x"6e207479",
  1330 => x"7065210d",
  1331 => x"00000000",
  1332 => x"436c7573",
  1333 => x"74657220",
  1334 => x"73697a65",
  1335 => x"3a202564",
  1336 => x"2c20436c",
  1337 => x"75737465",
  1338 => x"72206d61",
  1339 => x"736b2c20",
  1340 => x"25640a00",
  1341 => x"4f70656e",
  1342 => x"65642066",
  1343 => x"696c652c",
  1344 => x"206c6f61",
  1345 => x"64696e67",
  1346 => x"2e2e2e0a",
  1347 => x"00000000",
  1348 => x"43616e27",
  1349 => x"74206f70",
  1350 => x"656e2025",
  1351 => x"730a0000",
	others => x"00000000"
);

begin

process (clk)
begin
	if (clk'event and clk = '1') then
		if (from_zpu.memAWriteEnable = '1') and (from_zpu.memBWriteEnable = '1') and (from_zpu.memAAddr=from_zpu.memBAddr) and (from_zpu.memAWrite/=from_zpu.memBWrite) then
			report "write collision" severity failure;
		end if;
	
		if (from_zpu.memAWriteEnable = '1') then
			ram(to_integer(unsigned(from_zpu.memAAddr(maxAddrBitBRAM downto 2)))) := from_zpu.memAWrite;
			to_zpu.memARead <= from_zpu.memAWrite;
		else
			to_zpu.memARead <= ram(to_integer(unsigned(from_zpu.memAAddr(maxAddrBitBRAM downto 2))));
		end if;
	end if;
end process;

process (clk)
begin
	if (clk'event and clk = '1') then
		if (from_zpu.memBWriteEnable = '1') then
			ram(to_integer(unsigned(from_zpu.memBAddr(maxAddrBitBRAM downto 2)))) := from_zpu.memBWrite;
			to_zpu.memBRead <= from_zpu.memBWrite;
		else
			to_zpu.memBRead <= ram(to_integer(unsigned(from_zpu.memBAddr(maxAddrBitBRAM downto 2))));
		end if;
	end if;
end process;


end arch;

