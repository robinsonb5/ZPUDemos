-- ZPU
--
-- Copyright 2004-2008 oharboe - �yvind Harboe - oyvind.harboe@zylin.com
-- Modified by Alastair M. Robinson for the ZPUFlex project.
--
-- The FreeBSD license
-- 
-- Redistribution and use in source and binary forms, with or without
-- modification, are permitted provided that the following conditions
-- are met:
-- 
-- 1. Redistributions of source code must retain the above copyright
--    notice, this list of conditions and the following disclaimer.
-- 2. Redistributions in binary form must reproduce the above
--    copyright notice, this list of conditions and the following
--    disclaimer in the documentation and/or other materials
--    provided with the distribution.
-- 
-- THIS SOFTWARE IS PROVIDED BY THE ZPU PROJECT ``AS IS'' AND ANY
-- EXPRESS OR IMPLIED WARRANTIES, INCLUDING, BUT NOT LIMITED TO,
-- THE IMPLIED WARRANTIES OF MERCHANTABILITY AND FITNESS FOR A
-- PARTICULAR PURPOSE ARE DISCLAIMED. IN NO EVENT SHALL THE
-- ZPU PROJECT OR CONTRIBUTORS BE LIABLE FOR ANY DIRECT,
-- INDIRECT, INCIDENTAL, SPECIAL, EXEMPLARY, OR CONSEQUENTIAL DAMAGES
-- (INCLUDING, BUT NOT LIMITED TO, PROCUREMENT OF SUBSTITUTE GOODS
-- OR SERVICES; LOSS OF USE, DATA, OR PROFITS; OR BUSINESS INTERRUPTION)
-- HOWEVER CAUSED AND ON ANY THEORY OF LIABILITY, WHETHER IN CONTRACT,
-- STRICT LIABILITY, OR TORT (INCLUDING NEGLIGENCE OR OTHERWISE)
-- ARISING IN ANY WAY OUT OF THE USE OF THIS SOFTWARE, EVEN IF
-- ADVISED OF THE POSSIBILITY OF SUCH DAMAGE.
-- 
-- The views and conclusions contained in the software and documentation
-- are those of the authors and should not be interpreted as representing
-- official policies, either expressed or implied, of the ZPU Project.

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;


library work;
use work.zpupkg.all;

entity SDRAMTest_ROM is
generic
	(
		maxAddrBitBRAM : integer := maxAddrBitBRAMLimit -- Specify your actual ROM size to save LEs and unnecessary block RAM usage.
	);
port (
	clk : in std_logic;
	areset : in std_logic := '0';
	from_zpu : in ZPU_ToROM;
	to_zpu : out ZPU_FromROM
);
end SDRAMTest_ROM;

architecture arch of SDRAMTest_ROM is

type ram_type is array(natural range 0 to ((2**(maxAddrBitBRAM+1))/4)-1) of std_logic_vector(wordSize-1 downto 0);

shared variable ram : ram_type :=
(
     0 => x"84808080",
     1 => x"8c0b8480",
     2 => x"8081e004",
     3 => x"00848080",
     4 => x"808c04ff",
     5 => x"0d800404",
     6 => x"40000017",
     7 => x"00000000",
     8 => x"84808097",
     9 => x"fc088480",
    10 => x"80988008",
    11 => x"84808098",
    12 => x"84088480",
    13 => x"80809808",
    14 => x"2d848080",
    15 => x"98840c84",
    16 => x"80809880",
    17 => x"0c848080",
    18 => x"97fc0c04",
    19 => x"00000000",
    20 => x"00000000",
    21 => x"00000000",
    22 => x"00000000",
    23 => x"00000000",
    24 => x"71fd0608",
    25 => x"72830609",
    26 => x"81058205",
    27 => x"832b2a83",
    28 => x"ffff0652",
    29 => x"0471fc06",
    30 => x"08728306",
    31 => x"09810583",
    32 => x"05101010",
    33 => x"2a81ff06",
    34 => x"520471fd",
    35 => x"060883ff",
    36 => x"ff738306",
    37 => x"09810582",
    38 => x"05832b2b",
    39 => x"09067383",
    40 => x"ffff0673",
    41 => x"83060981",
    42 => x"05820583",
    43 => x"2b0b2b07",
    44 => x"72fc060c",
    45 => x"51510471",
    46 => x"fc060884",
    47 => x"808091f0",
    48 => x"73830610",
    49 => x"10050806",
    50 => x"7381ff06",
    51 => x"73830609",
    52 => x"81058305",
    53 => x"1010102b",
    54 => x"0772fc06",
    55 => x"0c515104",
    56 => x"84808097",
    57 => x"fc708480",
    58 => x"80999c27",
    59 => x"8e388071",
    60 => x"70840553",
    61 => x"0c848080",
    62 => x"81e50484",
    63 => x"8080808c",
    64 => x"51848080",
    65 => x"8edb0402",
    66 => x"c0050d02",
    67 => x"80c4055b",
    68 => x"80707c70",
    69 => x"84055e08",
    70 => x"725f5f5f",
    71 => x"5a7c7084",
    72 => x"055e0857",
    73 => x"80597698",
    74 => x"2a77882b",
    75 => x"58557480",
    76 => x"2e82f338",
    77 => x"7b802e80",
    78 => x"d338805c",
    79 => x"7480e42e",
    80 => x"81de3874",
    81 => x"80f82e81",
    82 => x"d7387480",
    83 => x"e42e81e2",
    84 => x"387480e4",
    85 => x"2680f138",
    86 => x"7480e32e",
    87 => x"80c838a5",
    88 => x"51848080",
    89 => x"868b2d74",
    90 => x"51848080",
    91 => x"868b2d82",
    92 => x"1a811a5a",
    93 => x"5a837925",
    94 => x"ffac3874",
    95 => x"ff9f387e",
    96 => x"84808097",
    97 => x"fc0c0280",
    98 => x"c0050d04",
    99 => x"74a52e09",
   100 => x"81069b38",
   101 => x"810b811a",
   102 => x"5a5c8379",
   103 => x"25ff8738",
   104 => x"84808082",
   105 => x"fb047a84",
   106 => x"1c710857",
   107 => x"5c547451",
   108 => x"84808086",
   109 => x"8b2d811a",
   110 => x"811a5a5a",
   111 => x"837925fe",
   112 => x"e5388480",
   113 => x"8082fb04",
   114 => x"7480f32e",
   115 => x"81e53874",
   116 => x"80f82e09",
   117 => x"8106ff87",
   118 => x"387d5380",
   119 => x"58777e24",
   120 => x"82963872",
   121 => x"802e81f9",
   122 => x"38875672",
   123 => x"9c2a7384",
   124 => x"2b545271",
   125 => x"802e8338",
   126 => x"8158b712",
   127 => x"54718924",
   128 => x"8438b012",
   129 => x"547780f0",
   130 => x"38ff1656",
   131 => x"758025db",
   132 => x"38811959",
   133 => x"837925fe",
   134 => x"8d388480",
   135 => x"8082fb04",
   136 => x"7a841c71",
   137 => x"08405c52",
   138 => x"7480e42e",
   139 => x"098106fe",
   140 => x"a0387d54",
   141 => x"8058777e",
   142 => x"24819538",
   143 => x"73802e81",
   144 => x"a0388756",
   145 => x"739c2a74",
   146 => x"842b5552",
   147 => x"71802e83",
   148 => x"388158b7",
   149 => x"12537189",
   150 => x"248438b0",
   151 => x"125377af",
   152 => x"38ff1656",
   153 => x"758025dc",
   154 => x"38811959",
   155 => x"837925fd",
   156 => x"b5388480",
   157 => x"8082fb04",
   158 => x"73518480",
   159 => x"80868b2d",
   160 => x"ff165675",
   161 => x"8025fee3",
   162 => x"38848080",
   163 => x"84910472",
   164 => x"51848080",
   165 => x"868b2dff",
   166 => x"16567580",
   167 => x"25ffa538",
   168 => x"84808084",
   169 => x"e9047984",
   170 => x"808097fc",
   171 => x"0c0280c0",
   172 => x"050d047a",
   173 => x"841c7108",
   174 => x"535c5384",
   175 => x"808086b0",
   176 => x"2d811959",
   177 => x"837925fc",
   178 => x"dd388480",
   179 => x"8082fb04",
   180 => x"ad518480",
   181 => x"80868b2d",
   182 => x"7d098105",
   183 => x"5473fee2",
   184 => x"38b05184",
   185 => x"8080868b",
   186 => x"2d811959",
   187 => x"837925fc",
   188 => x"b5388480",
   189 => x"8082fb04",
   190 => x"ad518480",
   191 => x"80868b2d",
   192 => x"7d098105",
   193 => x"53848080",
   194 => x"83e30402",
   195 => x"f8050d73",
   196 => x"52c00870",
   197 => x"882a7081",
   198 => x"06515151",
   199 => x"70802ef1",
   200 => x"3871c00c",
   201 => x"71848080",
   202 => x"97fc0c02",
   203 => x"88050d04",
   204 => x"02e8050d",
   205 => x"80785755",
   206 => x"75708405",
   207 => x"57085380",
   208 => x"5472982a",
   209 => x"73882b54",
   210 => x"5271802e",
   211 => x"a238c008",
   212 => x"70882a70",
   213 => x"81065151",
   214 => x"5170802e",
   215 => x"f13871c0",
   216 => x"0c811581",
   217 => x"15555583",
   218 => x"7425d638",
   219 => x"71ca3874",
   220 => x"84808097",
   221 => x"fc0c0298",
   222 => x"050d0402",
   223 => x"f4050d74",
   224 => x"76525380",
   225 => x"71259038",
   226 => x"70527270",
   227 => x"84055408",
   228 => x"ff135351",
   229 => x"71f43802",
   230 => x"8c050d04",
   231 => x"02d4050d",
   232 => x"7c7e5c58",
   233 => x"810b8480",
   234 => x"80928058",
   235 => x"5a835976",
   236 => x"08780c77",
   237 => x"08770856",
   238 => x"5473752e",
   239 => x"94387708",
   240 => x"53745284",
   241 => x"80809290",
   242 => x"51848080",
   243 => x"82872d80",
   244 => x"5a775680",
   245 => x"7b259038",
   246 => x"7a557570",
   247 => x"84055708",
   248 => x"ff165654",
   249 => x"74f43877",
   250 => x"08770856",
   251 => x"5675752e",
   252 => x"94387708",
   253 => x"53745284",
   254 => x"808092d0",
   255 => x"51848080",
   256 => x"82872d80",
   257 => x"5aff1984",
   258 => x"18585978",
   259 => x"8025ff9f",
   260 => x"38798480",
   261 => x"8097fc0c",
   262 => x"02ac050d",
   263 => x"0402e405",
   264 => x"0d787a55",
   265 => x"56815785",
   266 => x"aad5aad5",
   267 => x"760cfad5",
   268 => x"aad5aa0b",
   269 => x"8c170ccc",
   270 => x"7634b30b",
   271 => x"8f173475",
   272 => x"085372fc",
   273 => x"e2d5aad5",
   274 => x"2e923875",
   275 => x"08528480",
   276 => x"80939051",
   277 => x"84808082",
   278 => x"872d8057",
   279 => x"8c160855",
   280 => x"74fad5aa",
   281 => x"d4b32e93",
   282 => x"388c1608",
   283 => x"52848080",
   284 => x"93cc5184",
   285 => x"80808287",
   286 => x"2d805775",
   287 => x"55807425",
   288 => x"8e387470",
   289 => x"84055608",
   290 => x"ff155553",
   291 => x"73f43875",
   292 => x"085473fc",
   293 => x"e2d5aad5",
   294 => x"2e923875",
   295 => x"08528480",
   296 => x"80948851",
   297 => x"84808082",
   298 => x"872d8057",
   299 => x"8c160853",
   300 => x"72fad5aa",
   301 => x"d4b32e93",
   302 => x"388c1608",
   303 => x"52848080",
   304 => x"94c45184",
   305 => x"80808287",
   306 => x"2d805776",
   307 => x"84808097",
   308 => x"fc0c029c",
   309 => x"050d0402",
   310 => x"c4050d60",
   311 => x"5b806290",
   312 => x"808029ff",
   313 => x"05848080",
   314 => x"95805340",
   315 => x"5a848080",
   316 => x"82872d80",
   317 => x"e1b35780",
   318 => x"fe5eae51",
   319 => x"84808086",
   320 => x"8b2d7610",
   321 => x"70962a81",
   322 => x"06565774",
   323 => x"802e8538",
   324 => x"76810757",
   325 => x"76952a81",
   326 => x"06587780",
   327 => x"2e853876",
   328 => x"81325778",
   329 => x"77077f06",
   330 => x"775e598f",
   331 => x"ffff5876",
   332 => x"bfffff06",
   333 => x"707a3282",
   334 => x"2b7c1151",
   335 => x"57760c76",
   336 => x"1070962a",
   337 => x"81065657",
   338 => x"74802e85",
   339 => x"38768107",
   340 => x"5776952a",
   341 => x"81065574",
   342 => x"802e8538",
   343 => x"76813257",
   344 => x"ff185877",
   345 => x"8025c838",
   346 => x"7c578fff",
   347 => x"ff5876bf",
   348 => x"ffff0670",
   349 => x"7a32822b",
   350 => x"7c057008",
   351 => x"575e5674",
   352 => x"762e80ea",
   353 => x"38807a53",
   354 => x"84808095",
   355 => x"90525c84",
   356 => x"80808287",
   357 => x"2d745475",
   358 => x"53755284",
   359 => x"808095a4",
   360 => x"51848080",
   361 => x"82872d7b",
   362 => x"5a761070",
   363 => x"962a8106",
   364 => x"57577580",
   365 => x"2e853876",
   366 => x"81075776",
   367 => x"952a8106",
   368 => x"5574802e",
   369 => x"85387681",
   370 => x"3257ff18",
   371 => x"58778025",
   372 => x"ff9c38ff",
   373 => x"1e5e7dfe",
   374 => x"a1388a51",
   375 => x"84808086",
   376 => x"8b2d7b84",
   377 => x"808097fc",
   378 => x"0c02bc05",
   379 => x"0d04811a",
   380 => x"5a848080",
   381 => x"8ba90402",
   382 => x"cc050d7e",
   383 => x"605e5881",
   384 => x"5a805b80",
   385 => x"c07a585c",
   386 => x"85ada989",
   387 => x"bb780c79",
   388 => x"59815697",
   389 => x"55767607",
   390 => x"822b7811",
   391 => x"515485ad",
   392 => x"a989bb74",
   393 => x"0c7510ff",
   394 => x"16565674",
   395 => x"8025e638",
   396 => x"7610811a",
   397 => x"5a579879",
   398 => x"25d73877",
   399 => x"56807d25",
   400 => x"90387c55",
   401 => x"75708405",
   402 => x"5708ff16",
   403 => x"565474f4",
   404 => x"388157ff",
   405 => x"8787a5c3",
   406 => x"780c9759",
   407 => x"76822b78",
   408 => x"1170085f",
   409 => x"56567cff",
   410 => x"8787a5c3",
   411 => x"2e80cc38",
   412 => x"74085473",
   413 => x"85ada989",
   414 => x"bb2e9438",
   415 => x"80750854",
   416 => x"76538480",
   417 => x"8095cc52",
   418 => x"5a848080",
   419 => x"82872d76",
   420 => x"10ff1a5a",
   421 => x"57788025",
   422 => x"c3387a82",
   423 => x"2b5675b1",
   424 => x"387b5284",
   425 => x"808095ec",
   426 => x"51848080",
   427 => x"82872d7b",
   428 => x"84808097",
   429 => x"fc0c02b4",
   430 => x"050d047a",
   431 => x"77077710",
   432 => x"ff1b5b58",
   433 => x"5b788025",
   434 => x"ff923884",
   435 => x"80808d9a",
   436 => x"04755284",
   437 => x"808096a8",
   438 => x"51848080",
   439 => x"82872d75",
   440 => x"992a8132",
   441 => x"81067009",
   442 => x"81057107",
   443 => x"7009709f",
   444 => x"2c7d0679",
   445 => x"109fffff",
   446 => x"fc066081",
   447 => x"2a415a5d",
   448 => x"57585975",
   449 => x"da387909",
   450 => x"8105707b",
   451 => x"079f2a55",
   452 => x"567bbf26",
   453 => x"8438739d",
   454 => x"38817053",
   455 => x"84808095",
   456 => x"ec525c84",
   457 => x"80808287",
   458 => x"2d7b8480",
   459 => x"8097fc0c",
   460 => x"02b4050d",
   461 => x"04848080",
   462 => x"96c05184",
   463 => x"80808287",
   464 => x"2d7b5284",
   465 => x"808095ec",
   466 => x"51848080",
   467 => x"82872d7b",
   468 => x"84808097",
   469 => x"fc0c02b4",
   470 => x"050d0402",
   471 => x"dc050d81",
   472 => x"0b848080",
   473 => x"92805858",
   474 => x"83597608",
   475 => x"800c8008",
   476 => x"77085654",
   477 => x"73752e94",
   478 => x"38800853",
   479 => x"74528480",
   480 => x"80929051",
   481 => x"84808082",
   482 => x"872d8058",
   483 => x"80705755",
   484 => x"75708405",
   485 => x"57088116",
   486 => x"5654a080",
   487 => x"7524f138",
   488 => x"80087708",
   489 => x"56567575",
   490 => x"2e943880",
   491 => x"08537452",
   492 => x"84808092",
   493 => x"d0518480",
   494 => x"8082872d",
   495 => x"8058ff19",
   496 => x"84185859",
   497 => x"788025ff",
   498 => x"a1387780",
   499 => x"2e8d3884",
   500 => x"8080978c",
   501 => x"51848080",
   502 => x"82872d81",
   503 => x"5785aad5",
   504 => x"aad50b80",
   505 => x"0cfad5aa",
   506 => x"d5aa0b8c",
   507 => x"0ccc0b80",
   508 => x"34b30b8f",
   509 => x"34800855",
   510 => x"74fce2d5",
   511 => x"aad52e92",
   512 => x"38800852",
   513 => x"84808093",
   514 => x"90518480",
   515 => x"8082872d",
   516 => x"80578c08",
   517 => x"5877fad5",
   518 => x"aad4b32e",
   519 => x"92388c08",
   520 => x"52848080",
   521 => x"93cc5184",
   522 => x"80808287",
   523 => x"2d805780",
   524 => x"70575575",
   525 => x"70840557",
   526 => x"08811656",
   527 => x"54a08075",
   528 => x"24f13880",
   529 => x"085978fc",
   530 => x"e2d5aad5",
   531 => x"2e923880",
   532 => x"08528480",
   533 => x"80948851",
   534 => x"84808082",
   535 => x"872d8057",
   536 => x"8c085473",
   537 => x"fad5aad4",
   538 => x"b32e80ea",
   539 => x"388c0852",
   540 => x"84808094",
   541 => x"c4518480",
   542 => x"8082872d",
   543 => x"a0805280",
   544 => x"51848080",
   545 => x"8bf72d84",
   546 => x"808097fc",
   547 => x"08548480",
   548 => x"8097fc08",
   549 => x"802e8d38",
   550 => x"84808097",
   551 => x"b0518480",
   552 => x"8082872d",
   553 => x"73528051",
   554 => x"84808089",
   555 => x"d72d8480",
   556 => x"8097fc08",
   557 => x"802efda7",
   558 => x"38848080",
   559 => x"97c85184",
   560 => x"80808287",
   561 => x"2d810b84",
   562 => x"80809280",
   563 => x"58588359",
   564 => x"8480808e",
   565 => x"ea047680",
   566 => x"2effa138",
   567 => x"84808097",
   568 => x"e0518480",
   569 => x"8082872d",
   570 => x"84808090",
   571 => x"fc040000",
   572 => x"00ffffff",
   573 => x"ff00ffff",
   574 => x"ffff00ff",
   575 => x"ffffff00",
   576 => x"00000000",
   577 => x"55555555",
   578 => x"aaaaaaaa",
   579 => x"ffffffff",
   580 => x"53616e69",
   581 => x"74792063",
   582 => x"6865636b",
   583 => x"20666169",
   584 => x"6c656420",
   585 => x"28626566",
   586 => x"6f726520",
   587 => x"63616368",
   588 => x"65207265",
   589 => x"66726573",
   590 => x"6829206f",
   591 => x"6e203078",
   592 => x"25642028",
   593 => x"676f7420",
   594 => x"30782564",
   595 => x"290a0000",
   596 => x"53616e69",
   597 => x"74792063",
   598 => x"6865636b",
   599 => x"20666169",
   600 => x"6c656420",
   601 => x"28616674",
   602 => x"65722063",
   603 => x"61636865",
   604 => x"20726566",
   605 => x"72657368",
   606 => x"29206f6e",
   607 => x"20307825",
   608 => x"64202867",
   609 => x"6f742030",
   610 => x"78256429",
   611 => x"0a000000",
   612 => x"42797465",
   613 => x"20636865",
   614 => x"636b2066",
   615 => x"61696c65",
   616 => x"64202862",
   617 => x"65666f72",
   618 => x"65206361",
   619 => x"63686520",
   620 => x"72656672",
   621 => x"65736829",
   622 => x"20617420",
   623 => x"30202867",
   624 => x"6f742030",
   625 => x"78256429",
   626 => x"0a000000",
   627 => x"42797465",
   628 => x"20636865",
   629 => x"636b2066",
   630 => x"61696c65",
   631 => x"64202862",
   632 => x"65666f72",
   633 => x"65206361",
   634 => x"63686520",
   635 => x"72656672",
   636 => x"65736829",
   637 => x"20617420",
   638 => x"33202867",
   639 => x"6f742030",
   640 => x"78256429",
   641 => x"0a000000",
   642 => x"42797465",
   643 => x"20636865",
   644 => x"636b2066",
   645 => x"61696c65",
   646 => x"64202861",
   647 => x"66746572",
   648 => x"20636163",
   649 => x"68652072",
   650 => x"65667265",
   651 => x"73682920",
   652 => x"61742030",
   653 => x"2028676f",
   654 => x"74203078",
   655 => x"2564290a",
   656 => x"00000000",
   657 => x"42797465",
   658 => x"20636865",
   659 => x"636b2066",
   660 => x"61696c65",
   661 => x"64202861",
   662 => x"66746572",
   663 => x"20636163",
   664 => x"68652072",
   665 => x"65667265",
   666 => x"73682920",
   667 => x"61742033",
   668 => x"2028676f",
   669 => x"74203078",
   670 => x"2564290a",
   671 => x"00000000",
   672 => x"43686563",
   673 => x"6b696e67",
   674 => x"206d656d",
   675 => x"6f727900",
   676 => x"30782564",
   677 => x"20676f6f",
   678 => x"64207265",
   679 => x"6164732c",
   680 => x"20000000",
   681 => x"4572726f",
   682 => x"72206174",
   683 => x"20307825",
   684 => x"642c2065",
   685 => x"78706563",
   686 => x"74656420",
   687 => x"30782564",
   688 => x"2c20676f",
   689 => x"74203078",
   690 => x"25640a00",
   691 => x"42616420",
   692 => x"64617461",
   693 => x"20666f75",
   694 => x"6e642061",
   695 => x"74203078",
   696 => x"25642028",
   697 => x"30782564",
   698 => x"290a0000",
   699 => x"53445241",
   700 => x"4d207369",
   701 => x"7a652028",
   702 => x"61737375",
   703 => x"6d696e67",
   704 => x"206e6f20",
   705 => x"61646472",
   706 => x"65737320",
   707 => x"6661756c",
   708 => x"74732920",
   709 => x"69732030",
   710 => x"78256420",
   711 => x"6d656761",
   712 => x"62797465",
   713 => x"730a0000",
   714 => x"416c6961",
   715 => x"73657320",
   716 => x"666f756e",
   717 => x"64206174",
   718 => x"20307825",
   719 => x"640a0000",
   720 => x"28416c69",
   721 => x"61736573",
   722 => x"2070726f",
   723 => x"6261626c",
   724 => x"79207369",
   725 => x"6d706c79",
   726 => x"20696e64",
   727 => x"69636174",
   728 => x"65207468",
   729 => x"61742052",
   730 => x"414d0a69",
   731 => x"7320736d",
   732 => x"616c6c65",
   733 => x"72207468",
   734 => x"616e2036",
   735 => x"34206d65",
   736 => x"67616279",
   737 => x"74657329",
   738 => x"0a000000",
   739 => x"46697273",
   740 => x"74207374",
   741 => x"61676520",
   742 => x"73616e69",
   743 => x"74792063",
   744 => x"6865636b",
   745 => x"20706173",
   746 => x"7365642e",
   747 => x"0a000000",
   748 => x"41646472",
   749 => x"65737320",
   750 => x"63686563",
   751 => x"6b207061",
   752 => x"73736564",
   753 => x"2e0a0000",
   754 => x"4c465352",
   755 => x"20636865",
   756 => x"636b2070",
   757 => x"61737365",
   758 => x"642e0a0a",
   759 => x"00000000",
   760 => x"42797465",
   761 => x"20286471",
   762 => x"6d292063",
   763 => x"6865636b",
   764 => x"20706173",
   765 => x"7365640a",
   766 => x"00000000",
	others => x"00000000"
);

begin

process (clk)
begin
	if (clk'event and clk = '1') then
		if (from_zpu.memAWriteEnable = '1') and (from_zpu.memBWriteEnable = '1') and (from_zpu.memAAddr=from_zpu.memBAddr) and (from_zpu.memAWrite/=from_zpu.memBWrite) then
			report "write collision" severity failure;
		end if;
	
		if (from_zpu.memAWriteEnable = '1') then
			ram(to_integer(unsigned(from_zpu.memAAddr(maxAddrBitBRAM downto 2)))) := from_zpu.memAWrite;
			to_zpu.memARead <= from_zpu.memAWrite;
		else
			to_zpu.memARead <= ram(to_integer(unsigned(from_zpu.memAAddr(maxAddrBitBRAM downto 2))));
		end if;
	end if;
end process;

process (clk)
begin
	if (clk'event and clk = '1') then
		if (from_zpu.memBWriteEnable = '1') then
			ram(to_integer(unsigned(from_zpu.memBAddr(maxAddrBitBRAM downto 2)))) := from_zpu.memBWrite;
			to_zpu.memBRead <= from_zpu.memBWrite;
		else
			to_zpu.memBRead <= ram(to_integer(unsigned(from_zpu.memBAddr(maxAddrBitBRAM downto 2))));
		end if;
	end if;
end process;


end arch;

