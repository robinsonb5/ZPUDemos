-- ZPU
--
-- Copyright 2004-2008 oharboe - �yvind Harboe - oyvind.harboe@zylin.com
-- Modified by Alastair M. Robinson for the ZPUFlex project.
--
-- The FreeBSD license
-- 
-- Redistribution and use in source and binary forms, with or without
-- modification, are permitted provided that the following conditions
-- are met:
-- 
-- 1. Redistributions of source code must retain the above copyright
--    notice, this list of conditions and the following disclaimer.
-- 2. Redistributions in binary form must reproduce the above
--    copyright notice, this list of conditions and the following
--    disclaimer in the documentation and/or other materials
--    provided with the distribution.
-- 
-- THIS SOFTWARE IS PROVIDED BY THE ZPU PROJECT ``AS IS'' AND ANY
-- EXPRESS OR IMPLIED WARRANTIES, INCLUDING, BUT NOT LIMITED TO,
-- THE IMPLIED WARRANTIES OF MERCHANTABILITY AND FITNESS FOR A
-- PARTICULAR PURPOSE ARE DISCLAIMED. IN NO EVENT SHALL THE
-- ZPU PROJECT OR CONTRIBUTORS BE LIABLE FOR ANY DIRECT,
-- INDIRECT, INCIDENTAL, SPECIAL, EXEMPLARY, OR CONSEQUENTIAL DAMAGES
-- (INCLUDING, BUT NOT LIMITED TO, PROCUREMENT OF SUBSTITUTE GOODS
-- OR SERVICES; LOSS OF USE, DATA, OR PROFITS; OR BUSINESS INTERRUPTION)
-- HOWEVER CAUSED AND ON ANY THEORY OF LIABILITY, WHETHER IN CONTRACT,
-- STRICT LIABILITY, OR TORT (INCLUDING NEGLIGENCE OR OTHERWISE)
-- ARISING IN ANY WAY OUT OF THE USE OF THIS SOFTWARE, EVEN IF
-- ADVISED OF THE POSSIBILITY OF SUCH DAMAGE.
-- 
-- The views and conclusions contained in the software and documentation
-- are those of the authors and should not be interpreted as representing
-- official policies, either expressed or implied, of the ZPU Project.

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;


library work;
use work.zpu_config.all;
use work.zpupkg.all;

entity SDBootstrap_ROM is
generic
	(
		maxAddrBit : integer := maxAddrBitBRAMLimit -- Specify your actual ROM size to save LEs and unnecessary block RAM usage.
	);
port (
	clk : in std_logic;
	areset : in std_logic := '0';
	from_zpu : in ZPU_ToROM;
	to_zpu : out ZPU_FromROM
);
end SDBootstrap_ROM;

architecture arch of SDBootstrap_ROM is

type ram_type is array(natural range 0 to ((2**(maxAddrBit+1))/4)-1) of std_logic_vector(wordSize-1 downto 0);

shared variable ram : ram_type :=
(
     0 => x"0ba08080",
     1 => x"ec040000",
     2 => x"00000000",
     3 => x"0ba08080",
     4 => x"880d8004",
     5 => x"a0808094",
     6 => x"0471fd06",
     7 => x"08728306",
     8 => x"09810582",
     9 => x"05832b2a",
    10 => x"83ffff06",
    11 => x"520471fc",
    12 => x"06087283",
    13 => x"06098105",
    14 => x"83051010",
    15 => x"102a81ff",
    16 => x"06520471",
    17 => x"fc06080b",
    18 => x"a0809ee8",
    19 => x"73830610",
    20 => x"10050806",
    21 => x"7381ff06",
    22 => x"73830609",
    23 => x"81058305",
    24 => x"1010102b",
    25 => x"0772fc06",
    26 => x"0c515104",
    27 => x"0284050b",
    28 => x"a0808088",
    29 => x"0ca08080",
    30 => x"940ba080",
    31 => x"8d9b0400",
    32 => x"0002c405",
    33 => x"0d0280c0",
    34 => x"0583ffe0",
    35 => x"e05b5680",
    36 => x"76708405",
    37 => x"5808715e",
    38 => x"5e577c70",
    39 => x"84055e08",
    40 => x"58805b77",
    41 => x"982a7888",
    42 => x"2b595372",
    43 => x"8838765e",
    44 => x"a08083aa",
    45 => x"047b802e",
    46 => x"81ca3880",
    47 => x"5c7280e4",
    48 => x"2e9f3872",
    49 => x"80e4268d",
    50 => x"387280e3",
    51 => x"2e80ee38",
    52 => x"a08082ca",
    53 => x"047280f3",
    54 => x"2e80cc38",
    55 => x"a08082ca",
    56 => x"04758417",
    57 => x"71087e5c",
    58 => x"56575287",
    59 => x"55739c2a",
    60 => x"74842b55",
    61 => x"5271802e",
    62 => x"83388159",
    63 => x"89722589",
    64 => x"38b71252",
    65 => x"a080828c",
    66 => x"04b01252",
    67 => x"78802e88",
    68 => x"387151a0",
    69 => x"8083b52d",
    70 => x"ff155574",
    71 => x"8025ce38",
    72 => x"8054a080",
    73 => x"82e00475",
    74 => x"84177108",
    75 => x"70545c57",
    76 => x"52a08083",
    77 => x"d92d7b54",
    78 => x"a08082e0",
    79 => x"04758417",
    80 => x"71085557",
    81 => x"52a08083",
    82 => x"9304a551",
    83 => x"a08083b5",
    84 => x"2d7251a0",
    85 => x"8083b52d",
    86 => x"821757a0",
    87 => x"80839d04",
    88 => x"73ff1555",
    89 => x"52807225",
    90 => x"b4387970",
    91 => x"81055ba0",
    92 => x"8080ae2d",
    93 => x"705253a0",
    94 => x"8083b52d",
    95 => x"811757a0",
    96 => x"8082e004",
    97 => x"72a52e09",
    98 => x"81068838",
    99 => x"815ca080",
   100 => x"839d0472",
   101 => x"51a08083",
   102 => x"b52d8117",
   103 => x"57811b5b",
   104 => x"837b25fd",
   105 => x"fe3872fd",
   106 => x"f1387d83",
   107 => x"ffe0800c",
   108 => x"02bc050d",
   109 => x"0402f805",
   110 => x"0d7352c0",
   111 => x"0870882a",
   112 => x"70810651",
   113 => x"51517080",
   114 => x"2ef13871",
   115 => x"c00c7183",
   116 => x"ffe0800c",
   117 => x"0288050d",
   118 => x"0402e805",
   119 => x"0d775574",
   120 => x"70840556",
   121 => x"08538054",
   122 => x"72982a73",
   123 => x"882b5452",
   124 => x"71802ea2",
   125 => x"38c00870",
   126 => x"882a7081",
   127 => x"06515151",
   128 => x"70802ef1",
   129 => x"3871c00c",
   130 => x"81168115",
   131 => x"55568374",
   132 => x"25d63871",
   133 => x"ca387583",
   134 => x"ffe0800c",
   135 => x"0298050d",
   136 => x"0402f405",
   137 => x"0d747671",
   138 => x"81ff06d4",
   139 => x"0c535383",
   140 => x"fff1a008",
   141 => x"85387189",
   142 => x"2b527198",
   143 => x"2ad40c71",
   144 => x"902a7081",
   145 => x"ff06d40c",
   146 => x"5171882a",
   147 => x"7081ff06",
   148 => x"d40c5171",
   149 => x"81ff06d4",
   150 => x"0c72902a",
   151 => x"7081ff06",
   152 => x"d40c51d4",
   153 => x"087081ff",
   154 => x"06515182",
   155 => x"b8bf5270",
   156 => x"81ff2e09",
   157 => x"81069438",
   158 => x"81ff0bd4",
   159 => x"0cd40870",
   160 => x"81ff06ff",
   161 => x"14545151",
   162 => x"71e53870",
   163 => x"83ffe080",
   164 => x"0c028c05",
   165 => x"0d0402fc",
   166 => x"050d81c7",
   167 => x"5181ff0b",
   168 => x"d40cff11",
   169 => x"51708025",
   170 => x"f4380284",
   171 => x"050d0402",
   172 => x"f0050da0",
   173 => x"8085962d",
   174 => x"819c9f53",
   175 => x"805287fc",
   176 => x"80f751a0",
   177 => x"8084a12d",
   178 => x"83ffe080",
   179 => x"085483ff",
   180 => x"e0800881",
   181 => x"2e098106",
   182 => x"ab3881ff",
   183 => x"0bd40c82",
   184 => x"0a52849c",
   185 => x"80e951a0",
   186 => x"8084a12d",
   187 => x"83ffe080",
   188 => x"088d3881",
   189 => x"ff0bd40c",
   190 => x"7353a080",
   191 => x"868b04a0",
   192 => x"8085962d",
   193 => x"ff135372",
   194 => x"ffb23872",
   195 => x"83ffe080",
   196 => x"0c029005",
   197 => x"0d0402f4",
   198 => x"050d81ff",
   199 => x"0bd40ca0",
   200 => x"809ef851",
   201 => x"a08083d9",
   202 => x"2d935380",
   203 => x"5287fc80",
   204 => x"c151a080",
   205 => x"84a12d83",
   206 => x"ffe08008",
   207 => x"8d3881ff",
   208 => x"0bd40c81",
   209 => x"53a08086",
   210 => x"d504a080",
   211 => x"85962dff",
   212 => x"135372d7",
   213 => x"387283ff",
   214 => x"e0800c02",
   215 => x"8c050d04",
   216 => x"02f0050d",
   217 => x"a0808596",
   218 => x"2d83aa52",
   219 => x"849c80c8",
   220 => x"51a08084",
   221 => x"a12d83ff",
   222 => x"e0800883",
   223 => x"ffe08008",
   224 => x"53a0809f",
   225 => x"845254a0",
   226 => x"8081812d",
   227 => x"73812e09",
   228 => x"81069038",
   229 => x"d8087083",
   230 => x"ffff0654",
   231 => x"547283aa",
   232 => x"2ea338a0",
   233 => x"8086962d",
   234 => x"a08087be",
   235 => x"048154a0",
   236 => x"8088f304",
   237 => x"a0809f9c",
   238 => x"51a08081",
   239 => x"812d8054",
   240 => x"a08088f3",
   241 => x"047352a0",
   242 => x"809fb851",
   243 => x"a0808181",
   244 => x"2d81ff0b",
   245 => x"d40cb153",
   246 => x"a08085af",
   247 => x"2d83ffe0",
   248 => x"8008802e",
   249 => x"80f43880",
   250 => x"5287fc80",
   251 => x"fa51a080",
   252 => x"84a12d83",
   253 => x"ffe08008",
   254 => x"80d03883",
   255 => x"ffe08008",
   256 => x"52a0809f",
   257 => x"d051a080",
   258 => x"81812d81",
   259 => x"ff0bd40c",
   260 => x"d40881ff",
   261 => x"067053a0",
   262 => x"809fdc52",
   263 => x"54a08081",
   264 => x"812d81ff",
   265 => x"0bd40c81",
   266 => x"ff0bd40c",
   267 => x"81ff0bd4",
   268 => x"0c81ff0b",
   269 => x"d40c7386",
   270 => x"2a708106",
   271 => x"70565153",
   272 => x"72802eaf",
   273 => x"38a08087",
   274 => x"ad0483ff",
   275 => x"e0800852",
   276 => x"a0809fd0",
   277 => x"51a08081",
   278 => x"812d7282",
   279 => x"2efed538",
   280 => x"ff135372",
   281 => x"fef238a0",
   282 => x"809fec51",
   283 => x"a08083d9",
   284 => x"2d725473",
   285 => x"83ffe080",
   286 => x"0c029005",
   287 => x"0d0402f4",
   288 => x"050d810b",
   289 => x"83fff1a0",
   290 => x"0cd00870",
   291 => x"8f2a7081",
   292 => x"06515153",
   293 => x"72f33872",
   294 => x"d00ca080",
   295 => x"85962da0",
   296 => x"80a08451",
   297 => x"a08083d9",
   298 => x"2dd00870",
   299 => x"8f2a7081",
   300 => x"06515153",
   301 => x"72f33881",
   302 => x"0bd00c87",
   303 => x"53805284",
   304 => x"d480c051",
   305 => x"a08084a1",
   306 => x"2d83ffe0",
   307 => x"8008812e",
   308 => x"09810687",
   309 => x"3883ffe0",
   310 => x"800853a0",
   311 => x"80a09451",
   312 => x"a08083d9",
   313 => x"2d72822e",
   314 => x"09810692",
   315 => x"38a080a0",
   316 => x"a851a080",
   317 => x"83d92d80",
   318 => x"53a0808a",
   319 => x"ee04ff13",
   320 => x"5372ffb9",
   321 => x"38a080a0",
   322 => x"c851a080",
   323 => x"83d92da0",
   324 => x"8086e02d",
   325 => x"83ffe080",
   326 => x"0883fff1",
   327 => x"a00c83ff",
   328 => x"e0800880",
   329 => x"2e8b38a0",
   330 => x"80a0e451",
   331 => x"a08083d9",
   332 => x"2da080a0",
   333 => x"f851a080",
   334 => x"83d92d81",
   335 => x"5287fc80",
   336 => x"d051a080",
   337 => x"84a12d81",
   338 => x"ff0bd40c",
   339 => x"d008708f",
   340 => x"2a708106",
   341 => x"51515372",
   342 => x"f33872d0",
   343 => x"0c81ff0b",
   344 => x"d40ca080",
   345 => x"a18851a0",
   346 => x"8083d92d",
   347 => x"81537283",
   348 => x"ffe0800c",
   349 => x"028c050d",
   350 => x"04800b83",
   351 => x"ffe0800c",
   352 => x"0402e005",
   353 => x"0d797b57",
   354 => x"57805881",
   355 => x"ff0bd40c",
   356 => x"d008708f",
   357 => x"2a708106",
   358 => x"51515473",
   359 => x"f3388281",
   360 => x"0bd00c81",
   361 => x"ff0bd40c",
   362 => x"765287fc",
   363 => x"80d151a0",
   364 => x"8084a12d",
   365 => x"80dbc6df",
   366 => x"5583ffe0",
   367 => x"8008802e",
   368 => x"983883ff",
   369 => x"e0800853",
   370 => x"7652a080",
   371 => x"a19451a0",
   372 => x"8081812d",
   373 => x"a0808ca5",
   374 => x"0481ff0b",
   375 => x"d40cd408",
   376 => x"7081ff06",
   377 => x"51547381",
   378 => x"fe2e0981",
   379 => x"069b3880",
   380 => x"ff55d808",
   381 => x"76708405",
   382 => x"580cff15",
   383 => x"55748025",
   384 => x"f1388158",
   385 => x"a0808c8f",
   386 => x"04ff1555",
   387 => x"74cb3881",
   388 => x"ff0bd40c",
   389 => x"d008708f",
   390 => x"2a708106",
   391 => x"51515473",
   392 => x"f33873d0",
   393 => x"0c7783ff",
   394 => x"e0800c02",
   395 => x"a0050d04",
   396 => x"02f4050d",
   397 => x"7470882a",
   398 => x"83fe8006",
   399 => x"7072982a",
   400 => x"0772882b",
   401 => x"87fc8080",
   402 => x"0673982b",
   403 => x"81f00a06",
   404 => x"71730707",
   405 => x"83ffe080",
   406 => x"0c565153",
   407 => x"51028c05",
   408 => x"0d0402f8",
   409 => x"050d028e",
   410 => x"05a08080",
   411 => x"ae2d7498",
   412 => x"2b71902b",
   413 => x"0770902c",
   414 => x"83ffe080",
   415 => x"0c525202",
   416 => x"88050d04",
   417 => x"02f8050d",
   418 => x"7370902b",
   419 => x"71902a07",
   420 => x"83ffe080",
   421 => x"0c520288",
   422 => x"050d0402",
   423 => x"ec050d80",
   424 => x"0b870a0c",
   425 => x"a080a1b4",
   426 => x"51a08083",
   427 => x"d92da080",
   428 => x"88fe2d83",
   429 => x"ffe08008",
   430 => x"802e81e6",
   431 => x"38a080a1",
   432 => x"cc51a080",
   433 => x"83d92da0",
   434 => x"8090802d",
   435 => x"83ffe1a0",
   436 => x"52a080a1",
   437 => x"e451a080",
   438 => x"9c892d83",
   439 => x"ffe08008",
   440 => x"802e81be",
   441 => x"3883ffe1",
   442 => x"a00ba080",
   443 => x"a1f05254",
   444 => x"a08083d9",
   445 => x"2d805573",
   446 => x"70810555",
   447 => x"a08080ae",
   448 => x"2d5372a0",
   449 => x"2e80de38",
   450 => x"72a32e80",
   451 => x"fd387280",
   452 => x"c72e0981",
   453 => x"068b38a0",
   454 => x"80808c2d",
   455 => x"a0808ec1",
   456 => x"04728a2e",
   457 => x"0981068b",
   458 => x"38a08080",
   459 => x"942da080",
   460 => x"8ec10472",
   461 => x"80cc2e09",
   462 => x"81068638",
   463 => x"83ffe1a0",
   464 => x"547281df",
   465 => x"06f00570",
   466 => x"81ff0651",
   467 => x"53b87327",
   468 => x"8938ef13",
   469 => x"7081ff06",
   470 => x"51537484",
   471 => x"2b730755",
   472 => x"a0808df7",
   473 => x"0472a32e",
   474 => x"a1387370",
   475 => x"810555a0",
   476 => x"8080ae2d",
   477 => x"5372a02e",
   478 => x"f138ff14",
   479 => x"75537052",
   480 => x"54a0809c",
   481 => x"892d7487",
   482 => x"0a0c7370",
   483 => x"810555a0",
   484 => x"8080ae2d",
   485 => x"53728a2e",
   486 => x"098106ee",
   487 => x"38a0808d",
   488 => x"f504a080",
   489 => x"a28451a0",
   490 => x"8083d92d",
   491 => x"800b83ff",
   492 => x"e0800c02",
   493 => x"94050d04",
   494 => x"02e8050d",
   495 => x"77797b58",
   496 => x"55558053",
   497 => x"727625ab",
   498 => x"38747081",
   499 => x"0556a080",
   500 => x"80ae2d74",
   501 => x"70810556",
   502 => x"a08080ae",
   503 => x"2d525271",
   504 => x"712e8838",
   505 => x"8151a080",
   506 => x"8ff50481",
   507 => x"1353a080",
   508 => x"8fc40480",
   509 => x"517083ff",
   510 => x"e0800c02",
   511 => x"98050d04",
   512 => x"02d8050d",
   513 => x"ff0b83ff",
   514 => x"f5cc0c80",
   515 => x"0b83fff5",
   516 => x"e00ca080",
   517 => x"a29051a0",
   518 => x"8083d92d",
   519 => x"83fff1b8",
   520 => x"528051a0",
   521 => x"808b812d",
   522 => x"83ffe080",
   523 => x"085483ff",
   524 => x"e0800892",
   525 => x"38a080a2",
   526 => x"a051a080",
   527 => x"83d92d73",
   528 => x"55a08097",
   529 => x"e404a080",
   530 => x"a2b451a0",
   531 => x"8083d92d",
   532 => x"8056810b",
   533 => x"83fff1ac",
   534 => x"0c8853a0",
   535 => x"80a2cc52",
   536 => x"83fff1ee",
   537 => x"51a0808f",
   538 => x"b82d83ff",
   539 => x"e0800876",
   540 => x"2e098106",
   541 => x"8b3883ff",
   542 => x"e0800883",
   543 => x"fff1ac0c",
   544 => x"8853a080",
   545 => x"a2d85283",
   546 => x"fff28a51",
   547 => x"a0808fb8",
   548 => x"2d83ffe0",
   549 => x"80088b38",
   550 => x"83ffe080",
   551 => x"0883fff1",
   552 => x"ac0c83ff",
   553 => x"f1ac0852",
   554 => x"a080a2e4",
   555 => x"51a08081",
   556 => x"812d83ff",
   557 => x"f1ac0880",
   558 => x"2e81bb38",
   559 => x"83fff4fe",
   560 => x"0ba08080",
   561 => x"ae2d83ff",
   562 => x"f4ff0ba0",
   563 => x"8080ae2d",
   564 => x"71982b71",
   565 => x"902b0783",
   566 => x"fff5800b",
   567 => x"a08080ae",
   568 => x"2d70882b",
   569 => x"720783ff",
   570 => x"f5810ba0",
   571 => x"8080ae2d",
   572 => x"710783ff",
   573 => x"f5b60ba0",
   574 => x"8080ae2d",
   575 => x"83fff5b7",
   576 => x"0ba08080",
   577 => x"ae2d7188",
   578 => x"2b07535f",
   579 => x"54525a56",
   580 => x"57557381",
   581 => x"abaa2e09",
   582 => x"81069338",
   583 => x"7551a080",
   584 => x"8cb02d83",
   585 => x"ffe08008",
   586 => x"56a08092",
   587 => x"c4047382",
   588 => x"d4d52e90",
   589 => x"38a080a2",
   590 => x"f851a080",
   591 => x"83d92da0",
   592 => x"8094bc04",
   593 => x"7552a080",
   594 => x"a39851a0",
   595 => x"8081812d",
   596 => x"83fff1b8",
   597 => x"527551a0",
   598 => x"808b812d",
   599 => x"83ffe080",
   600 => x"085583ff",
   601 => x"e0800880",
   602 => x"2e84f938",
   603 => x"a080a3b0",
   604 => x"51a08083",
   605 => x"d92da080",
   606 => x"a3d851a0",
   607 => x"8081812d",
   608 => x"8853a080",
   609 => x"a2d85283",
   610 => x"fff28a51",
   611 => x"a0808fb8",
   612 => x"2d83ffe0",
   613 => x"80088d38",
   614 => x"810b83ff",
   615 => x"f5e00ca0",
   616 => x"8093cd04",
   617 => x"8853a080",
   618 => x"a2cc5283",
   619 => x"fff1ee51",
   620 => x"a0808fb8",
   621 => x"2d83ffe0",
   622 => x"8008802e",
   623 => x"9038a080",
   624 => x"a3f051a0",
   625 => x"8081812d",
   626 => x"a08094bc",
   627 => x"0483fff5",
   628 => x"b60ba080",
   629 => x"80ae2d54",
   630 => x"7380d52e",
   631 => x"09810680",
   632 => x"db3883ff",
   633 => x"f5b70ba0",
   634 => x"8080ae2d",
   635 => x"547381aa",
   636 => x"2e098106",
   637 => x"80c63880",
   638 => x"0b83fff1",
   639 => x"b80ba080",
   640 => x"80ae2d56",
   641 => x"547481e9",
   642 => x"2e833881",
   643 => x"547481eb",
   644 => x"2e8c3880",
   645 => x"5573752e",
   646 => x"09810683",
   647 => x"c73883ff",
   648 => x"f1c30ba0",
   649 => x"8080ae2d",
   650 => x"55749138",
   651 => x"83fff1c4",
   652 => x"0ba08080",
   653 => x"ae2d5473",
   654 => x"822e8838",
   655 => x"8055a080",
   656 => x"97e40483",
   657 => x"fff1c50b",
   658 => x"a08080ae",
   659 => x"2d7083ff",
   660 => x"f5e80cff",
   661 => x"0583fff5",
   662 => x"dc0c83ff",
   663 => x"f1c60ba0",
   664 => x"8080ae2d",
   665 => x"83fff1c7",
   666 => x"0ba08080",
   667 => x"ae2d5876",
   668 => x"05778280",
   669 => x"29057083",
   670 => x"fff5d00c",
   671 => x"83fff1c8",
   672 => x"0ba08080",
   673 => x"ae2d7083",
   674 => x"fff5c80c",
   675 => x"83fff5e0",
   676 => x"08595758",
   677 => x"76802e81",
   678 => x"df388853",
   679 => x"a080a2d8",
   680 => x"5283fff2",
   681 => x"8a51a080",
   682 => x"8fb82d83",
   683 => x"ffe08008",
   684 => x"82b23883",
   685 => x"fff5e808",
   686 => x"70842b83",
   687 => x"fff5b80c",
   688 => x"7083fff5",
   689 => x"e40c83ff",
   690 => x"f1dd0ba0",
   691 => x"8080ae2d",
   692 => x"83fff1dc",
   693 => x"0ba08080",
   694 => x"ae2d7182",
   695 => x"80290583",
   696 => x"fff1de0b",
   697 => x"a08080ae",
   698 => x"2d708480",
   699 => x"80291283",
   700 => x"fff1df0b",
   701 => x"a08080ae",
   702 => x"2d708180",
   703 => x"0a291270",
   704 => x"83fff1b0",
   705 => x"0c83fff5",
   706 => x"c8087129",
   707 => x"83fff5d0",
   708 => x"08057083",
   709 => x"fff5f00c",
   710 => x"83fff1e5",
   711 => x"0ba08080",
   712 => x"ae2d83ff",
   713 => x"f1e40ba0",
   714 => x"8080ae2d",
   715 => x"71828029",
   716 => x"0583fff1",
   717 => x"e60ba080",
   718 => x"80ae2d70",
   719 => x"84808029",
   720 => x"1283fff1",
   721 => x"e70ba080",
   722 => x"80ae2d70",
   723 => x"982b81f0",
   724 => x"0a067205",
   725 => x"7083fff1",
   726 => x"b40cfe11",
   727 => x"7e297705",
   728 => x"83fff5d8",
   729 => x"0c525952",
   730 => x"43545e51",
   731 => x"5259525d",
   732 => x"575957a0",
   733 => x"8097e204",
   734 => x"83fff1ca",
   735 => x"0ba08080",
   736 => x"ae2d83ff",
   737 => x"f1c90ba0",
   738 => x"8080ae2d",
   739 => x"71828029",
   740 => x"057083ff",
   741 => x"f5b80c70",
   742 => x"a02983ff",
   743 => x"0570892a",
   744 => x"7083fff5",
   745 => x"e40c83ff",
   746 => x"f1cf0ba0",
   747 => x"8080ae2d",
   748 => x"83fff1ce",
   749 => x"0ba08080",
   750 => x"ae2d7182",
   751 => x"80290570",
   752 => x"83fff1b0",
   753 => x"0c7b7129",
   754 => x"1e7083ff",
   755 => x"f5d80c7d",
   756 => x"83fff1b4",
   757 => x"0c730583",
   758 => x"fff5f00c",
   759 => x"555e5151",
   760 => x"55558155",
   761 => x"7483ffe0",
   762 => x"800c02a8",
   763 => x"050d0402",
   764 => x"ec050d76",
   765 => x"70872c71",
   766 => x"80ff0657",
   767 => x"555383ff",
   768 => x"f5e0088a",
   769 => x"3872882c",
   770 => x"7381ff06",
   771 => x"56547383",
   772 => x"fff5cc08",
   773 => x"2ea83883",
   774 => x"fff1b852",
   775 => x"83fff5d0",
   776 => x"081451a0",
   777 => x"808b812d",
   778 => x"83ffe080",
   779 => x"085383ff",
   780 => x"e0800880",
   781 => x"2e80cb38",
   782 => x"7383fff5",
   783 => x"cc0c83ff",
   784 => x"f5e00880",
   785 => x"2ea03874",
   786 => x"842983ff",
   787 => x"f1b80570",
   788 => x"085253a0",
   789 => x"808cb02d",
   790 => x"83ffe080",
   791 => x"08f00a06",
   792 => x"55a08099",
   793 => x"80047410",
   794 => x"83fff1b8",
   795 => x"0570a080",
   796 => x"80992d52",
   797 => x"53a0808c",
   798 => x"e22d83ff",
   799 => x"e0800855",
   800 => x"74537283",
   801 => x"ffe0800c",
   802 => x"0294050d",
   803 => x"0402cc05",
   804 => x"0d7e605e",
   805 => x"5b8056ff",
   806 => x"0b83fff5",
   807 => x"cc0c83ff",
   808 => x"f1b40883",
   809 => x"fff5d808",
   810 => x"565783ff",
   811 => x"f5e00876",
   812 => x"2e8e3883",
   813 => x"fff5e808",
   814 => x"842b59a0",
   815 => x"8099c804",
   816 => x"83fff5e4",
   817 => x"08842b59",
   818 => x"805a7979",
   819 => x"2781e138",
   820 => x"798f06a0",
   821 => x"17575473",
   822 => x"a1387452",
   823 => x"a080a490",
   824 => x"51a08081",
   825 => x"812d83ff",
   826 => x"f1b85274",
   827 => x"51811555",
   828 => x"a0808b81",
   829 => x"2d83fff1",
   830 => x"b8568076",
   831 => x"a08080ae",
   832 => x"2d555873",
   833 => x"782e8338",
   834 => x"81587381",
   835 => x"e52e8198",
   836 => x"38817079",
   837 => x"06555c73",
   838 => x"802e818c",
   839 => x"388b16a0",
   840 => x"8080ae2d",
   841 => x"98065877",
   842 => x"80fe388b",
   843 => x"537c5275",
   844 => x"51a0808f",
   845 => x"b82d83ff",
   846 => x"e0800880",
   847 => x"eb389c16",
   848 => x"0851a080",
   849 => x"8cb02d83",
   850 => x"ffe08008",
   851 => x"841c0c9a",
   852 => x"16a08080",
   853 => x"992d51a0",
   854 => x"808ce22d",
   855 => x"83ffe080",
   856 => x"0883ffe0",
   857 => x"80085555",
   858 => x"83fff5e0",
   859 => x"08802e9e",
   860 => x"389416a0",
   861 => x"8080992d",
   862 => x"51a0808c",
   863 => x"e22d83ff",
   864 => x"e0800890",
   865 => x"2b83fff0",
   866 => x"0a067016",
   867 => x"51547388",
   868 => x"1c0c777b",
   869 => x"0c7c52a0",
   870 => x"80a4b051",
   871 => x"a0808181",
   872 => x"2d7b54a0",
   873 => x"809bfe04",
   874 => x"811a5aa0",
   875 => x"8099ca04",
   876 => x"83fff5e0",
   877 => x"08802e80",
   878 => x"c3387651",
   879 => x"a08097ef",
   880 => x"2d83ffe0",
   881 => x"800883ff",
   882 => x"e0800853",
   883 => x"a080a4c4",
   884 => x"5257a080",
   885 => x"81812d76",
   886 => x"80ffffff",
   887 => x"f8065473",
   888 => x"80ffffff",
   889 => x"f82e9538",
   890 => x"fe1783ff",
   891 => x"f5e80829",
   892 => x"83fff5f0",
   893 => x"080555a0",
   894 => x"8099c804",
   895 => x"80547383",
   896 => x"ffe0800c",
   897 => x"02b4050d",
   898 => x"0402e405",
   899 => x"0d787a71",
   900 => x"5483fff5",
   901 => x"bc535555",
   902 => x"a080998d",
   903 => x"2d83ffe0",
   904 => x"800881ff",
   905 => x"06537280",
   906 => x"2e818338",
   907 => x"a080a4dc",
   908 => x"51a08083",
   909 => x"d92d83ff",
   910 => x"f5c00883",
   911 => x"ff05892a",
   912 => x"57807056",
   913 => x"56757725",
   914 => x"81803883",
   915 => x"fff5c408",
   916 => x"fe0583ff",
   917 => x"f5e80829",
   918 => x"83fff5f0",
   919 => x"08117683",
   920 => x"fff5dc08",
   921 => x"06057554",
   922 => x"5253a080",
   923 => x"8b812d83",
   924 => x"ffe08008",
   925 => x"802e80c7",
   926 => x"38811570",
   927 => x"83fff5dc",
   928 => x"08065455",
   929 => x"72963883",
   930 => x"fff5c408",
   931 => x"51a08097",
   932 => x"ef2d83ff",
   933 => x"e0800883",
   934 => x"fff5c40c",
   935 => x"84801481",
   936 => x"17575476",
   937 => x"7624ffa3",
   938 => x"38a0809d",
   939 => x"ca047452",
   940 => x"a080a4f8",
   941 => x"51a08081",
   942 => x"812da080",
   943 => x"9dcc0483",
   944 => x"ffe08008",
   945 => x"53a0809d",
   946 => x"cc048153",
   947 => x"7283ffe0",
   948 => x"800c029c",
   949 => x"050d0483",
   950 => x"ffe08c08",
   951 => x"0283ffe0",
   952 => x"8c0cff3d",
   953 => x"0d800b83",
   954 => x"ffe08c08",
   955 => x"fc050c83",
   956 => x"ffe08c08",
   957 => x"88050881",
   958 => x"06ff1170",
   959 => x"097083ff",
   960 => x"e08c088c",
   961 => x"05080683",
   962 => x"ffe08c08",
   963 => x"fc050811",
   964 => x"83ffe08c",
   965 => x"08fc050c",
   966 => x"83ffe08c",
   967 => x"08880508",
   968 => x"812a83ff",
   969 => x"e08c0888",
   970 => x"050c83ff",
   971 => x"e08c088c",
   972 => x"05081083",
   973 => x"ffe08c08",
   974 => x"8c050c51",
   975 => x"51515183",
   976 => x"ffe08c08",
   977 => x"88050880",
   978 => x"2e8438ff",
   979 => x"a23983ff",
   980 => x"e08c08fc",
   981 => x"05087083",
   982 => x"ffe0800c",
   983 => x"51833d0d",
   984 => x"83ffe08c",
   985 => x"0c040000",
   986 => x"00ffffff",
   987 => x"ff00ffff",
   988 => x"ffff00ff",
   989 => x"ffffff00",
   990 => x"436d645f",
   991 => x"696e6974",
   992 => x"0a000000",
   993 => x"636d645f",
   994 => x"434d4438",
   995 => x"20726573",
   996 => x"706f6e73",
   997 => x"653a2025",
   998 => x"640a0000",
   999 => x"53444843",
  1000 => x"20496e69",
  1001 => x"7469616c",
  1002 => x"697a6174",
  1003 => x"696f6e20",
  1004 => x"6572726f",
  1005 => x"72210a00",
  1006 => x"434d4438",
  1007 => x"5f342072",
  1008 => x"6573706f",
  1009 => x"6e73653a",
  1010 => x"2025640a",
  1011 => x"00000000",
  1012 => x"434d4435",
  1013 => x"38202564",
  1014 => x"0a202000",
  1015 => x"434d4435",
  1016 => x"385f3220",
  1017 => x"25640a20",
  1018 => x"20000000",
  1019 => x"44657465",
  1020 => x"726d696e",
  1021 => x"65642053",
  1022 => x"44484320",
  1023 => x"73746174",
  1024 => x"75730a00",
  1025 => x"41637469",
  1026 => x"76617469",
  1027 => x"6e672043",
  1028 => x"530a0000",
  1029 => x"53656e74",
  1030 => x"20726573",
  1031 => x"65742063",
  1032 => x"6f6d6d61",
  1033 => x"6e640a00",
  1034 => x"53442063",
  1035 => x"61726420",
  1036 => x"696e6974",
  1037 => x"69616c69",
  1038 => x"7a617469",
  1039 => x"6f6e2065",
  1040 => x"72726f72",
  1041 => x"210a0000",
  1042 => x"43617264",
  1043 => x"20726573",
  1044 => x"706f6e64",
  1045 => x"65642074",
  1046 => x"6f207265",
  1047 => x"7365740a",
  1048 => x"00000000",
  1049 => x"53444843",
  1050 => x"20636172",
  1051 => x"64206465",
  1052 => x"74656374",
  1053 => x"65640a00",
  1054 => x"53656e64",
  1055 => x"696e6720",
  1056 => x"636d6431",
  1057 => x"360a0000",
  1058 => x"496e6974",
  1059 => x"20646f6e",
  1060 => x"650a0000",
  1061 => x"52656164",
  1062 => x"20636f6d",
  1063 => x"6d616e64",
  1064 => x"20666169",
  1065 => x"6c656420",
  1066 => x"61742025",
  1067 => x"64202825",
  1068 => x"64290a00",
  1069 => x"496e6974",
  1070 => x"69616c69",
  1071 => x"7a696e67",
  1072 => x"20534420",
  1073 => x"63617264",
  1074 => x"0a000000",
  1075 => x"48756e74",
  1076 => x"696e6720",
  1077 => x"666f7220",
  1078 => x"70617274",
  1079 => x"6974696f",
  1080 => x"6e0a0000",
  1081 => x"4d414e49",
  1082 => x"46455354",
  1083 => x"4d535400",
  1084 => x"50617273",
  1085 => x"696e6720",
  1086 => x"6d616e69",
  1087 => x"66657374",
  1088 => x"0a000000",
  1089 => x"52657475",
  1090 => x"726e696e",
  1091 => x"670a0000",
  1092 => x"52656164",
  1093 => x"696e6720",
  1094 => x"4d42520a",
  1095 => x"00000000",
  1096 => x"52656164",
  1097 => x"206f6620",
  1098 => x"4d425220",
  1099 => x"6661696c",
  1100 => x"65640a00",
  1101 => x"4d425220",
  1102 => x"73756363",
  1103 => x"65737366",
  1104 => x"756c6c79",
  1105 => x"20726561",
  1106 => x"640a0000",
  1107 => x"46415431",
  1108 => x"36202020",
  1109 => x"00000000",
  1110 => x"46415433",
  1111 => x"32202020",
  1112 => x"00000000",
  1113 => x"50617274",
  1114 => x"6974696f",
  1115 => x"6e636f75",
  1116 => x"6e742025",
  1117 => x"640a0000",
  1118 => x"4e6f2070",
  1119 => x"61727469",
  1120 => x"74696f6e",
  1121 => x"20736967",
  1122 => x"6e617475",
  1123 => x"72652066",
  1124 => x"6f756e64",
  1125 => x"0a000000",
  1126 => x"52656164",
  1127 => x"696e6720",
  1128 => x"626f6f74",
  1129 => x"20736563",
  1130 => x"746f7220",
  1131 => x"25640a00",
  1132 => x"52656164",
  1133 => x"20626f6f",
  1134 => x"74207365",
  1135 => x"63746f72",
  1136 => x"2066726f",
  1137 => x"6d206669",
  1138 => x"72737420",
  1139 => x"70617274",
  1140 => x"6974696f",
  1141 => x"6e0a0000",
  1142 => x"48756e74",
  1143 => x"696e6720",
  1144 => x"666f7220",
  1145 => x"66696c65",
  1146 => x"73797374",
  1147 => x"656d0a00",
  1148 => x"556e7375",
  1149 => x"70706f72",
  1150 => x"74656420",
  1151 => x"70617274",
  1152 => x"6974696f",
  1153 => x"6e207479",
  1154 => x"7065210d",
  1155 => x"00000000",
  1156 => x"52656164",
  1157 => x"696e6720",
  1158 => x"64697265",
  1159 => x"63746f72",
  1160 => x"79207365",
  1161 => x"63746f72",
  1162 => x"2025640a",
  1163 => x"00000000",
  1164 => x"66696c65",
  1165 => x"20222573",
  1166 => x"2220666f",
  1167 => x"756e640d",
  1168 => x"00000000",
  1169 => x"47657446",
  1170 => x"41544c69",
  1171 => x"6e6b2072",
  1172 => x"65747572",
  1173 => x"6e656420",
  1174 => x"25640a00",
  1175 => x"4f70656e",
  1176 => x"65642066",
  1177 => x"696c652c",
  1178 => x"206c6f61",
  1179 => x"64696e67",
  1180 => x"2e2e2e0a",
  1181 => x"00000000",
  1182 => x"43616e27",
  1183 => x"74206f70",
  1184 => x"656e2025",
  1185 => x"730a0000",
	others => x"00000000"
);

begin

process (clk)
begin
	if (clk'event and clk = '1') then
		if (from_zpu.memAWriteEnable = '1') and (from_zpu.memBWriteEnable = '1') and (from_zpu.memAAddr=from_zpu.memBAddr) and (from_zpu.memAWrite/=from_zpu.memBWrite) then
			report "write collision" severity failure;
		end if;
	
		if (from_zpu.memAWriteEnable = '1') then
			ram(to_integer(unsigned(from_zpu.memAAddr(maxAddrBit downto 2)))) := from_zpu.memAWrite;
			to_zpu.memARead <= from_zpu.memAWrite;
		else
			to_zpu.memARead <= ram(to_integer(unsigned(from_zpu.memAAddr(maxAddrBit downto 2))));
		end if;
	end if;
end process;

process (clk)
begin
	if (clk'event and clk = '1') then
		if (from_zpu.memBWriteEnable = '1') then
			ram(to_integer(unsigned(from_zpu.memBAddr(maxAddrBit downto 2)))) := from_zpu.memBWrite;
			to_zpu.memBRead <= from_zpu.memBWrite;
		else
			to_zpu.memBRead <= ram(to_integer(unsigned(from_zpu.memBAddr(maxAddrBit downto 2))));
		end if;
	end if;
end process;


end arch;

