-- ZPU
--
-- Copyright 2004-2008 oharboe - �yvind Harboe - oyvind.harboe@zylin.com
-- Modified by Alastair M. Robinson for the ZPUFlex project.
--
-- The FreeBSD license
-- 
-- Redistribution and use in source and binary forms, with or without
-- modification, are permitted provided that the following conditions
-- are met:
-- 
-- 1. Redistributions of source code must retain the above copyright
--    notice, this list of conditions and the following disclaimer.
-- 2. Redistributions in binary form must reproduce the above
--    copyright notice, this list of conditions and the following
--    disclaimer in the documentation and/or other materials
--    provided with the distribution.
-- 
-- THIS SOFTWARE IS PROVIDED BY THE ZPU PROJECT ``AS IS'' AND ANY
-- EXPRESS OR IMPLIED WARRANTIES, INCLUDING, BUT NOT LIMITED TO,
-- THE IMPLIED WARRANTIES OF MERCHANTABILITY AND FITNESS FOR A
-- PARTICULAR PURPOSE ARE DISCLAIMED. IN NO EVENT SHALL THE
-- ZPU PROJECT OR CONTRIBUTORS BE LIABLE FOR ANY DIRECT,
-- INDIRECT, INCIDENTAL, SPECIAL, EXEMPLARY, OR CONSEQUENTIAL DAMAGES
-- (INCLUDING, BUT NOT LIMITED TO, PROCUREMENT OF SUBSTITUTE GOODS
-- OR SERVICES; LOSS OF USE, DATA, OR PROFITS; OR BUSINESS INTERRUPTION)
-- HOWEVER CAUSED AND ON ANY THEORY OF LIABILITY, WHETHER IN CONTRACT,
-- STRICT LIABILITY, OR TORT (INCLUDING NEGLIGENCE OR OTHERWISE)
-- ARISING IN ANY WAY OUT OF THE USE OF THIS SOFTWARE, EVEN IF
-- ADVISED OF THE POSSIBILITY OF SUCH DAMAGE.
-- 
-- The views and conclusions contained in the software and documentation
-- are those of the authors and should not be interpreted as representing
-- official policies, either expressed or implied, of the ZPU Project.

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;


library work;
use work.zpu_config.all;
use work.zpupkg.all;

entity SDRAMTest_ROM is
generic
	(
		maxAddrBitBRAM : integer := maxAddrBitBRAMLimit -- Specify your actual ROM size to save LEs and unnecessary block RAM usage.
	);
port (
	clk : in std_logic;
	areset : in std_logic := '0';
	from_zpu : in ZPU_ToROM;
	to_zpu : out ZPU_FromROM
);
end SDRAMTest_ROM;

architecture arch of SDRAMTest_ROM is

type ram_type is array(natural range 0 to ((2**(maxAddrBitBRAM+1))/4)-1) of std_logic_vector(wordSize-1 downto 0);

shared variable ram : ram_type :=
(
     0 => x"0ba08080",
     1 => x"ec040000",
     2 => x"00000000",
     3 => x"0ba08080",
     4 => x"880d8004",
     5 => x"a0808094",
     6 => x"0471fd06",
     7 => x"08728306",
     8 => x"09810582",
     9 => x"05832b2a",
    10 => x"83ffff06",
    11 => x"520471fc",
    12 => x"06087283",
    13 => x"06098105",
    14 => x"83051010",
    15 => x"102a81ff",
    16 => x"06520471",
    17 => x"fc06080b",
    18 => x"a0808ee8",
    19 => x"73830610",
    20 => x"10050806",
    21 => x"7381ff06",
    22 => x"73830609",
    23 => x"81058305",
    24 => x"1010102b",
    25 => x"0772fc06",
    26 => x"0c515104",
    27 => x"0284050b",
    28 => x"a0808088",
    29 => x"0ca08080",
    30 => x"940ba080",
    31 => x"8bf20400",
    32 => x"0002c005",
    33 => x"0d0280c4",
    34 => x"05a08095",
    35 => x"d45c5c80",
    36 => x"7c708405",
    37 => x"5e08715f",
    38 => x"5f587d70",
    39 => x"84055f08",
    40 => x"57805a76",
    41 => x"982a7788",
    42 => x"2b585574",
    43 => x"802e8291",
    44 => x"387c802e",
    45 => x"80c23880",
    46 => x"5d7480e4",
    47 => x"2e81b238",
    48 => x"7480e426",
    49 => x"80eb3874",
    50 => x"80e32e80",
    51 => x"c438a551",
    52 => x"a08083cd",
    53 => x"2d7451a0",
    54 => x"8083cd2d",
    55 => x"82185881",
    56 => x"1a5a837a",
    57 => x"25ffbc38",
    58 => x"74ffaf38",
    59 => x"7ea08094",
    60 => x"f40c0280",
    61 => x"c0050d04",
    62 => x"74a52e09",
    63 => x"81069a38",
    64 => x"810b811b",
    65 => x"5b5d837a",
    66 => x"25ff9838",
    67 => x"a08081e8",
    68 => x"047b841d",
    69 => x"7108575d",
    70 => x"547451a0",
    71 => x"8083cd2d",
    72 => x"8118811b",
    73 => x"5b58837a",
    74 => x"25fef838",
    75 => x"a08081e8",
    76 => x"047480f3",
    77 => x"2e098106",
    78 => x"ff94387b",
    79 => x"841d7108",
    80 => x"70545d5d",
    81 => x"53a08083",
    82 => x"f12d800b",
    83 => x"ff115452",
    84 => x"807225ff",
    85 => x"8a387a70",
    86 => x"81055c33",
    87 => x"705255a0",
    88 => x"8083cd2d",
    89 => x"811873ff",
    90 => x"15555358",
    91 => x"a08082d0",
    92 => x"047b841d",
    93 => x"71087f5c",
    94 => x"555d5287",
    95 => x"56729c2a",
    96 => x"73842b54",
    97 => x"5271802e",
    98 => x"83388159",
    99 => x"b7125471",
   100 => x"89248438",
   101 => x"b0125478",
   102 => x"9438ff16",
   103 => x"56758025",
   104 => x"dc38800b",
   105 => x"ff115452",
   106 => x"a08082d0",
   107 => x"047351a0",
   108 => x"8083cd2d",
   109 => x"ff165675",
   110 => x"8025c238",
   111 => x"a08083a2",
   112 => x"0477a080",
   113 => x"94f40c02",
   114 => x"80c0050d",
   115 => x"0402f805",
   116 => x"0d7352c0",
   117 => x"0870882a",
   118 => x"70810651",
   119 => x"51517080",
   120 => x"2ef13871",
   121 => x"c00c71a0",
   122 => x"8094f40c",
   123 => x"0288050d",
   124 => x"0402e805",
   125 => x"0d807857",
   126 => x"55757084",
   127 => x"05570853",
   128 => x"80547298",
   129 => x"2a73882b",
   130 => x"54527180",
   131 => x"2ea238c0",
   132 => x"0870882a",
   133 => x"70810651",
   134 => x"51517080",
   135 => x"2ef13871",
   136 => x"c00c8115",
   137 => x"81155555",
   138 => x"837425d6",
   139 => x"3871ca38",
   140 => x"74a08094",
   141 => x"f40c0298",
   142 => x"050d0402",
   143 => x"f4050d74",
   144 => x"76525380",
   145 => x"71259038",
   146 => x"70527270",
   147 => x"84055408",
   148 => x"ff135351",
   149 => x"71f43802",
   150 => x"8c050d04",
   151 => x"02d4050d",
   152 => x"7c7e5c58",
   153 => x"810ba080",
   154 => x"8ef8585a",
   155 => x"83597608",
   156 => x"780c7708",
   157 => x"77085654",
   158 => x"73752e92",
   159 => x"38770853",
   160 => x"7452a080",
   161 => x"8f8851a0",
   162 => x"8081812d",
   163 => x"805a7756",
   164 => x"807b2590",
   165 => x"387a5575",
   166 => x"70840557",
   167 => x"08ff1656",
   168 => x"5474f438",
   169 => x"77087708",
   170 => x"56567575",
   171 => x"2e923877",
   172 => x"08537452",
   173 => x"a0808fc8",
   174 => x"51a08081",
   175 => x"812d805a",
   176 => x"ff198418",
   177 => x"58597880",
   178 => x"25ffa338",
   179 => x"79a08094",
   180 => x"f40c02ac",
   181 => x"050d0402",
   182 => x"e4050d78",
   183 => x"7a555681",
   184 => x"5785aad5",
   185 => x"aad5760c",
   186 => x"fad5aad5",
   187 => x"aa0b8c17",
   188 => x"0ccc7634",
   189 => x"b30b8f17",
   190 => x"34750853",
   191 => x"72fce2d5",
   192 => x"aad52e90",
   193 => x"38750852",
   194 => x"a0809088",
   195 => x"51a08081",
   196 => x"812d8057",
   197 => x"8c160855",
   198 => x"74fad5aa",
   199 => x"d4b32e91",
   200 => x"388c1608",
   201 => x"52a08090",
   202 => x"c451a080",
   203 => x"81812d80",
   204 => x"57755580",
   205 => x"74258e38",
   206 => x"74708405",
   207 => x"5608ff15",
   208 => x"555373f4",
   209 => x"38750854",
   210 => x"73fce2d5",
   211 => x"aad52e90",
   212 => x"38750852",
   213 => x"a0809180",
   214 => x"51a08081",
   215 => x"812d8057",
   216 => x"8c160853",
   217 => x"72fad5aa",
   218 => x"d4b32e91",
   219 => x"388c1608",
   220 => x"52a08091",
   221 => x"bc51a080",
   222 => x"81812d80",
   223 => x"5776a080",
   224 => x"94f40c02",
   225 => x"9c050d04",
   226 => x"02c4050d",
   227 => x"605b8062",
   228 => x"90808029",
   229 => x"ff05a080",
   230 => x"91f85340",
   231 => x"5aa08081",
   232 => x"812d80e1",
   233 => x"b35780fe",
   234 => x"5eae51a0",
   235 => x"8083cd2d",
   236 => x"76107096",
   237 => x"2a810656",
   238 => x"5774802e",
   239 => x"85387681",
   240 => x"07577695",
   241 => x"2a810658",
   242 => x"77802e85",
   243 => x"38768132",
   244 => x"57787707",
   245 => x"7f06775e",
   246 => x"598fffff",
   247 => x"5876bfff",
   248 => x"ff06707a",
   249 => x"32822b7c",
   250 => x"11515776",
   251 => x"0c761070",
   252 => x"962a8106",
   253 => x"56577480",
   254 => x"2e853876",
   255 => x"81075776",
   256 => x"952a8106",
   257 => x"5574802e",
   258 => x"85387681",
   259 => x"3257ff18",
   260 => x"58778025",
   261 => x"c8387c57",
   262 => x"8fffff58",
   263 => x"76bfffff",
   264 => x"06707a32",
   265 => x"822b7c05",
   266 => x"7008575e",
   267 => x"5674762e",
   268 => x"80e43880",
   269 => x"7a53a080",
   270 => x"9288525c",
   271 => x"a0808181",
   272 => x"2d745475",
   273 => x"537552a0",
   274 => x"80929c51",
   275 => x"a0808181",
   276 => x"2d7b5a76",
   277 => x"1070962a",
   278 => x"81065757",
   279 => x"75802e85",
   280 => x"38768107",
   281 => x"5776952a",
   282 => x"81065574",
   283 => x"802e8538",
   284 => x"76813257",
   285 => x"ff185877",
   286 => x"8025ffa0",
   287 => x"38ff1e5e",
   288 => x"7dfea638",
   289 => x"8a51a080",
   290 => x"83cd2d7b",
   291 => x"a08094f4",
   292 => x"0c02bc05",
   293 => x"0d04811a",
   294 => x"5aa08088",
   295 => x"d30402cc",
   296 => x"050d7e60",
   297 => x"5e58815a",
   298 => x"805b80c0",
   299 => x"7a585c85",
   300 => x"ada989bb",
   301 => x"780c7959",
   302 => x"81569755",
   303 => x"76760782",
   304 => x"2b781151",
   305 => x"5485ada9",
   306 => x"89bb740c",
   307 => x"7510ff16",
   308 => x"56567480",
   309 => x"25e63876",
   310 => x"10811a5a",
   311 => x"57987925",
   312 => x"d7387756",
   313 => x"807d2590",
   314 => x"387c5575",
   315 => x"70840557",
   316 => x"08ff1656",
   317 => x"5474f438",
   318 => x"8157ff87",
   319 => x"87a5c378",
   320 => x"0c975976",
   321 => x"822b7811",
   322 => x"70085f56",
   323 => x"567cff87",
   324 => x"87a5c32e",
   325 => x"80c73874",
   326 => x"08547385",
   327 => x"ada989bb",
   328 => x"2e923880",
   329 => x"75085476",
   330 => x"53a08092",
   331 => x"c4525aa0",
   332 => x"8081812d",
   333 => x"7610ff1a",
   334 => x"5a577880",
   335 => x"25c5387a",
   336 => x"822b5675",
   337 => x"ad387b52",
   338 => x"a08092e4",
   339 => x"51a08081",
   340 => x"812d7ba0",
   341 => x"8094f40c",
   342 => x"02b4050d",
   343 => x"047a7707",
   344 => x"7710ff1b",
   345 => x"5b585b78",
   346 => x"8025ff97",
   347 => x"38a0808a",
   348 => x"bf047552",
   349 => x"a08093a0",
   350 => x"51a08081",
   351 => x"812d7599",
   352 => x"2a813281",
   353 => x"06700981",
   354 => x"05710770",
   355 => x"09709f2c",
   356 => x"7d067910",
   357 => x"9ffffffc",
   358 => x"0660812a",
   359 => x"415a5d57",
   360 => x"585975da",
   361 => x"38790981",
   362 => x"05707b07",
   363 => x"9f2a5556",
   364 => x"7bbf2684",
   365 => x"38739a38",
   366 => x"817053a0",
   367 => x"8092e452",
   368 => x"5ca08081",
   369 => x"812d7ba0",
   370 => x"8094f40c",
   371 => x"02b4050d",
   372 => x"04a08093",
   373 => x"b851a080",
   374 => x"81812d7b",
   375 => x"52a08092",
   376 => x"e451a080",
   377 => x"81812d7b",
   378 => x"a08094f4",
   379 => x"0c02b405",
   380 => x"0d0402dc",
   381 => x"050d810b",
   382 => x"a0808ef8",
   383 => x"58588359",
   384 => x"7608800c",
   385 => x"80087708",
   386 => x"56547375",
   387 => x"2e923880",
   388 => x"08537452",
   389 => x"a0808f88",
   390 => x"51a08081",
   391 => x"812d8058",
   392 => x"80705755",
   393 => x"75708405",
   394 => x"57088116",
   395 => x"5654a080",
   396 => x"7524f138",
   397 => x"80087708",
   398 => x"56567575",
   399 => x"2e923880",
   400 => x"08537452",
   401 => x"a0808fc8",
   402 => x"51a08081",
   403 => x"812d8058",
   404 => x"ff198418",
   405 => x"58597880",
   406 => x"25ffa538",
   407 => x"77802e8b",
   408 => x"38a08094",
   409 => x"8451a080",
   410 => x"81812d81",
   411 => x"5785aad5",
   412 => x"aad50b80",
   413 => x"0cfad5aa",
   414 => x"d5aa0b8c",
   415 => x"0ccc0b80",
   416 => x"34b30b8f",
   417 => x"34800855",
   418 => x"74fce2d5",
   419 => x"aad52e90",
   420 => x"38800852",
   421 => x"a0809088",
   422 => x"51a08081",
   423 => x"812d8057",
   424 => x"8c085877",
   425 => x"fad5aad4",
   426 => x"b32e9038",
   427 => x"8c0852a0",
   428 => x"8090c451",
   429 => x"a0808181",
   430 => x"2d805780",
   431 => x"70575575",
   432 => x"70840557",
   433 => x"08811656",
   434 => x"54a08075",
   435 => x"24f13880",
   436 => x"085978fc",
   437 => x"e2d5aad5",
   438 => x"2e903880",
   439 => x"0852a080",
   440 => x"918051a0",
   441 => x"8081812d",
   442 => x"80578c08",
   443 => x"5473fad5",
   444 => x"aad4b32e",
   445 => x"80dd388c",
   446 => x"0852a080",
   447 => x"91bc51a0",
   448 => x"8081812d",
   449 => x"a0805280",
   450 => x"51a08089",
   451 => x"9e2da080",
   452 => x"94f40854",
   453 => x"a08094f4",
   454 => x"08802e8b",
   455 => x"38a08094",
   456 => x"a851a080",
   457 => x"81812d73",
   458 => x"528051a0",
   459 => x"8087882d",
   460 => x"a08094f4",
   461 => x"08802efd",
   462 => x"bd38a080",
   463 => x"94c051a0",
   464 => x"8081812d",
   465 => x"810ba080",
   466 => x"8ef85858",
   467 => x"8359a080",
   468 => x"8c800476",
   469 => x"802effac",
   470 => x"38a08094",
   471 => x"d851a080",
   472 => x"81812da0",
   473 => x"808e8404",
   474 => x"00ffffff",
   475 => x"ff00ffff",
   476 => x"ffff00ff",
   477 => x"ffffff00",
   478 => x"00000000",
   479 => x"55555555",
   480 => x"aaaaaaaa",
   481 => x"ffffffff",
   482 => x"53616e69",
   483 => x"74792063",
   484 => x"6865636b",
   485 => x"20666169",
   486 => x"6c656420",
   487 => x"28626566",
   488 => x"6f726520",
   489 => x"63616368",
   490 => x"65207265",
   491 => x"66726573",
   492 => x"6829206f",
   493 => x"6e203078",
   494 => x"25642028",
   495 => x"676f7420",
   496 => x"30782564",
   497 => x"290a0000",
   498 => x"53616e69",
   499 => x"74792063",
   500 => x"6865636b",
   501 => x"20666169",
   502 => x"6c656420",
   503 => x"28616674",
   504 => x"65722063",
   505 => x"61636865",
   506 => x"20726566",
   507 => x"72657368",
   508 => x"29206f6e",
   509 => x"20307825",
   510 => x"64202867",
   511 => x"6f742030",
   512 => x"78256429",
   513 => x"0a000000",
   514 => x"42797465",
   515 => x"20636865",
   516 => x"636b2066",
   517 => x"61696c65",
   518 => x"64202862",
   519 => x"65666f72",
   520 => x"65206361",
   521 => x"63686520",
   522 => x"72656672",
   523 => x"65736829",
   524 => x"20617420",
   525 => x"30202867",
   526 => x"6f742030",
   527 => x"78256429",
   528 => x"0a000000",
   529 => x"42797465",
   530 => x"20636865",
   531 => x"636b2066",
   532 => x"61696c65",
   533 => x"64202862",
   534 => x"65666f72",
   535 => x"65206361",
   536 => x"63686520",
   537 => x"72656672",
   538 => x"65736829",
   539 => x"20617420",
   540 => x"33202867",
   541 => x"6f742030",
   542 => x"78256429",
   543 => x"0a000000",
   544 => x"42797465",
   545 => x"20636865",
   546 => x"636b2066",
   547 => x"61696c65",
   548 => x"64202861",
   549 => x"66746572",
   550 => x"20636163",
   551 => x"68652072",
   552 => x"65667265",
   553 => x"73682920",
   554 => x"61742030",
   555 => x"2028676f",
   556 => x"74203078",
   557 => x"2564290a",
   558 => x"00000000",
   559 => x"42797465",
   560 => x"20636865",
   561 => x"636b2066",
   562 => x"61696c65",
   563 => x"64202861",
   564 => x"66746572",
   565 => x"20636163",
   566 => x"68652072",
   567 => x"65667265",
   568 => x"73682920",
   569 => x"61742033",
   570 => x"2028676f",
   571 => x"74203078",
   572 => x"2564290a",
   573 => x"00000000",
   574 => x"43686563",
   575 => x"6b696e67",
   576 => x"206d656d",
   577 => x"6f727900",
   578 => x"30782564",
   579 => x"20676f6f",
   580 => x"64207265",
   581 => x"6164732c",
   582 => x"20000000",
   583 => x"4572726f",
   584 => x"72206174",
   585 => x"20307825",
   586 => x"642c2065",
   587 => x"78706563",
   588 => x"74656420",
   589 => x"30782564",
   590 => x"2c20676f",
   591 => x"74203078",
   592 => x"25640a00",
   593 => x"42616420",
   594 => x"64617461",
   595 => x"20666f75",
   596 => x"6e642061",
   597 => x"74203078",
   598 => x"25642028",
   599 => x"30782564",
   600 => x"290a0000",
   601 => x"53445241",
   602 => x"4d207369",
   603 => x"7a652028",
   604 => x"61737375",
   605 => x"6d696e67",
   606 => x"206e6f20",
   607 => x"61646472",
   608 => x"65737320",
   609 => x"6661756c",
   610 => x"74732920",
   611 => x"69732030",
   612 => x"78256420",
   613 => x"6d656761",
   614 => x"62797465",
   615 => x"730a0000",
   616 => x"416c6961",
   617 => x"73657320",
   618 => x"666f756e",
   619 => x"64206174",
   620 => x"20307825",
   621 => x"640a0000",
   622 => x"28416c69",
   623 => x"61736573",
   624 => x"2070726f",
   625 => x"6261626c",
   626 => x"79207369",
   627 => x"6d706c79",
   628 => x"20696e64",
   629 => x"69636174",
   630 => x"65207468",
   631 => x"61742052",
   632 => x"414d0a69",
   633 => x"7320736d",
   634 => x"616c6c65",
   635 => x"72207468",
   636 => x"616e2036",
   637 => x"34206d65",
   638 => x"67616279",
   639 => x"74657329",
   640 => x"0a000000",
   641 => x"46697273",
   642 => x"74207374",
   643 => x"61676520",
   644 => x"73616e69",
   645 => x"74792063",
   646 => x"6865636b",
   647 => x"20706173",
   648 => x"7365642e",
   649 => x"0a000000",
   650 => x"41646472",
   651 => x"65737320",
   652 => x"63686563",
   653 => x"6b207061",
   654 => x"73736564",
   655 => x"2e0a0000",
   656 => x"4c465352",
   657 => x"20636865",
   658 => x"636b2070",
   659 => x"61737365",
   660 => x"642e0a0a",
   661 => x"00000000",
   662 => x"42797465",
   663 => x"20286471",
   664 => x"6d292063",
   665 => x"6865636b",
   666 => x"20706173",
   667 => x"7365640a",
   668 => x"00000000",
	others => x"00000000"
);

begin

process (clk)
begin
	if (clk'event and clk = '1') then
		if (from_zpu.memAWriteEnable = '1') and (from_zpu.memBWriteEnable = '1') and (from_zpu.memAAddr=from_zpu.memBAddr) and (from_zpu.memAWrite/=from_zpu.memBWrite) then
			report "write collision" severity failure;
		end if;
	
		if (from_zpu.memAWriteEnable = '1') then
			ram(to_integer(unsigned(from_zpu.memAAddr(maxAddrBitBRAM downto 2)))) := from_zpu.memAWrite;
			to_zpu.memARead <= from_zpu.memAWrite;
		else
			to_zpu.memARead <= ram(to_integer(unsigned(from_zpu.memAAddr(maxAddrBitBRAM downto 2))));
		end if;
	end if;
end process;

process (clk)
begin
	if (clk'event and clk = '1') then
		if (from_zpu.memBWriteEnable = '1') then
			ram(to_integer(unsigned(from_zpu.memBAddr(maxAddrBitBRAM downto 2)))) := from_zpu.memBWrite;
			to_zpu.memBRead <= from_zpu.memBWrite;
		else
			to_zpu.memBRead <= ram(to_integer(unsigned(from_zpu.memBAddr(maxAddrBitBRAM downto 2))));
		end if;
	end if;
end process;


end arch;

