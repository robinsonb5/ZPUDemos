-- ZPU
--
-- Copyright 2004-2008 oharboe - �yvind Harboe - oyvind.harboe@zylin.com
-- Modified by Alastair M. Robinson for the ZPUFlex project.
--
-- The FreeBSD license
-- 
-- Redistribution and use in source and binary forms, with or without
-- modification, are permitted provided that the following conditions
-- are met:
-- 
-- 1. Redistributions of source code must retain the above copyright
--    notice, this list of conditions and the following disclaimer.
-- 2. Redistributions in binary form must reproduce the above
--    copyright notice, this list of conditions and the following
--    disclaimer in the documentation and/or other materials
--    provided with the distribution.
-- 
-- THIS SOFTWARE IS PROVIDED BY THE ZPU PROJECT ``AS IS'' AND ANY
-- EXPRESS OR IMPLIED WARRANTIES, INCLUDING, BUT NOT LIMITED TO,
-- THE IMPLIED WARRANTIES OF MERCHANTABILITY AND FITNESS FOR A
-- PARTICULAR PURPOSE ARE DISCLAIMED. IN NO EVENT SHALL THE
-- ZPU PROJECT OR CONTRIBUTORS BE LIABLE FOR ANY DIRECT,
-- INDIRECT, INCIDENTAL, SPECIAL, EXEMPLARY, OR CONSEQUENTIAL DAMAGES
-- (INCLUDING, BUT NOT LIMITED TO, PROCUREMENT OF SUBSTITUTE GOODS
-- OR SERVICES; LOSS OF USE, DATA, OR PROFITS; OR BUSINESS INTERRUPTION)
-- HOWEVER CAUSED AND ON ANY THEORY OF LIABILITY, WHETHER IN CONTRACT,
-- STRICT LIABILITY, OR TORT (INCLUDING NEGLIGENCE OR OTHERWISE)
-- ARISING IN ANY WAY OUT OF THE USE OF THIS SOFTWARE, EVEN IF
-- ADVISED OF THE POSSIBILITY OF SUCH DAMAGE.
-- 
-- The views and conclusions contained in the software and documentation
-- are those of the authors and should not be interpreted as representing
-- official policies, either expressed or implied, of the ZPU Project.

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;


library work;
use work.zpu_config.all;
use work.zpupkg.all;

entity RS232Bootstrap_ROM is
generic
	(
		maxAddrBitBRAM : integer := maxAddrBitBRAMLimit -- Specify your actual ROM size to save LEs and unnecessary block RAM usage.
	);
port (
	clk : in std_logic;
	areset : in std_logic := '0';
	from_zpu : in ZPU_ToROM;
	to_zpu : out ZPU_FromROM
);
end RS232Bootstrap_ROM;

architecture arch of RS232Bootstrap_ROM is

type ram_type is array(natural range 0 to ((2**(maxAddrBitBRAM+1))/4)-1) of std_logic_vector(wordSize-1 downto 0);

shared variable ram : ram_type :=
(
     0 => x"84808080",
     1 => x"ed040000",
     2 => x"00000000",
     3 => x"84808080",
     4 => x"880d8004",
     5 => x"84808080",
     6 => x"940471fd",
     7 => x"06087283",
     8 => x"06098105",
     9 => x"8205832b",
    10 => x"2a83ffff",
    11 => x"06520471",
    12 => x"fc060872",
    13 => x"83060981",
    14 => x"05830510",
    15 => x"10102a81",
    16 => x"ff065204",
    17 => x"71fc0608",
    18 => x"84808086",
    19 => x"b4738306",
    20 => x"10100508",
    21 => x"067381ff",
    22 => x"06738306",
    23 => x"09810583",
    24 => x"05101010",
    25 => x"2b0772fc",
    26 => x"060c5151",
    27 => x"04028405",
    28 => x"84808080",
    29 => x"880c8480",
    30 => x"8080940b",
    31 => x"84808085",
    32 => x"e0040000",
    33 => x"02f8050d",
    34 => x"7352c008",
    35 => x"70882a70",
    36 => x"81065151",
    37 => x"5170802e",
    38 => x"f13871c0",
    39 => x"0c7183ff",
    40 => x"e0800c02",
    41 => x"88050d04",
    42 => x"02e8050d",
    43 => x"80785755",
    44 => x"75708405",
    45 => x"57085380",
    46 => x"5472982a",
    47 => x"73882b54",
    48 => x"5271802e",
    49 => x"a238c008",
    50 => x"70882a70",
    51 => x"81065151",
    52 => x"5170802e",
    53 => x"f13871c0",
    54 => x"0c811581",
    55 => x"15555583",
    56 => x"7425d638",
    57 => x"71ca3874",
    58 => x"83ffe080",
    59 => x"0c029805",
    60 => x"0d0402f8",
    61 => x"050dc008",
    62 => x"70892a70",
    63 => x"81065152",
    64 => x"5270802e",
    65 => x"f1387181",
    66 => x"ff0683ff",
    67 => x"e0800c02",
    68 => x"88050d04",
    69 => x"02fc050d",
    70 => x"7381df06",
    71 => x"c9055170",
    72 => x"80258438",
    73 => x"a7115172",
    74 => x"842b7107",
    75 => x"83ffe080",
    76 => x"0c028405",
    77 => x"0d0402f0",
    78 => x"050d0297",
    79 => x"05848080",
    80 => x"80af2d83",
    81 => x"ffe0a408",
    82 => x"810583ff",
    83 => x"e0a40c54",
    84 => x"7380d32e",
    85 => x"098106a3",
    86 => x"38800b83",
    87 => x"ffe0a40c",
    88 => x"800b83ff",
    89 => x"e0940c80",
    90 => x"0b83ffe0",
    91 => x"a80c800b",
    92 => x"83ffe090",
    93 => x"0c848080",
    94 => x"85db0483",
    95 => x"ffe0a408",
    96 => x"5271812e",
    97 => x"09810680",
    98 => x"c13883ff",
    99 => x"e0900874",
   100 => x"81df06c9",
   101 => x"05525270",
   102 => x"80258438",
   103 => x"a7115171",
   104 => x"842b7107",
   105 => x"7083ffe0",
   106 => x"900c7052",
   107 => x"52837225",
   108 => x"85388a72",
   109 => x"31517010",
   110 => x"820583ff",
   111 => x"e09c0c80",
   112 => x"f40bc00c",
   113 => x"84808085",
   114 => x"db047183",
   115 => x"24a63883",
   116 => x"ffe0a808",
   117 => x"7481df06",
   118 => x"c9055252",
   119 => x"70802584",
   120 => x"38a71151",
   121 => x"71842b71",
   122 => x"0783ffe0",
   123 => x"a80c8480",
   124 => x"8085db04",
   125 => x"83ffe09c",
   126 => x"08830551",
   127 => x"717124a6",
   128 => x"3883ffe0",
   129 => x"94087481",
   130 => x"df06c905",
   131 => x"52527080",
   132 => x"258438a7",
   133 => x"11517184",
   134 => x"2b710783",
   135 => x"ffe0940c",
   136 => x"84808085",
   137 => x"950483ff",
   138 => x"e09008ff",
   139 => x"11525370",
   140 => x"82268197",
   141 => x"3883ffe0",
   142 => x"a8081081",
   143 => x"05517171",
   144 => x"2480df38",
   145 => x"83ffe0a0",
   146 => x"087481df",
   147 => x"06c90552",
   148 => x"52708025",
   149 => x"8438a711",
   150 => x"5171842b",
   151 => x"71077083",
   152 => x"ffe0a00c",
   153 => x"83ffe098",
   154 => x"08ff0583",
   155 => x"ffe0980c",
   156 => x"5283ffe0",
   157 => x"98088025",
   158 => x"80e13883",
   159 => x"ffe09408",
   160 => x"51717184",
   161 => x"808080c4",
   162 => x"2d83ffe0",
   163 => x"94088105",
   164 => x"83ffe094",
   165 => x"0c810b83",
   166 => x"ffe0980c",
   167 => x"84808085",
   168 => x"db0483ff",
   169 => x"e09808b3",
   170 => x"3883ffe0",
   171 => x"a008842b",
   172 => x"7083ffe0",
   173 => x"a00c83ff",
   174 => x"e0940852",
   175 => x"52717184",
   176 => x"808080c4",
   177 => x"2d848080",
   178 => x"85db0486",
   179 => x"73258c38",
   180 => x"80c20bc0",
   181 => x"0c848080",
   182 => x"808c2d02",
   183 => x"90050d04",
   184 => x"02fc050d",
   185 => x"80d25184",
   186 => x"80808184",
   187 => x"2d80e551",
   188 => x"84808081",
   189 => x"842d80e1",
   190 => x"51848080",
   191 => x"81842d80",
   192 => x"e4518480",
   193 => x"8081842d",
   194 => x"80f95184",
   195 => x"80808184",
   196 => x"2d8a5184",
   197 => x"80808184",
   198 => x"2d848080",
   199 => x"81f22d83",
   200 => x"ffe08008",
   201 => x"81ff0651",
   202 => x"84808082",
   203 => x"b62d8480",
   204 => x"80869904",
   205 => x"00ffffff",
   206 => x"ff00ffff",
   207 => x"ffff00ff",
   208 => x"ffffff00",
	others => x"00000000"
);

begin

process (clk)
begin
	if (clk'event and clk = '1') then
		if (from_zpu.memAWriteEnable = '1') and (from_zpu.memBWriteEnable = '1') and (from_zpu.memAAddr=from_zpu.memBAddr) and (from_zpu.memAWrite/=from_zpu.memBWrite) then
			report "write collision" severity failure;
		end if;
	
		if (from_zpu.memAWriteEnable = '1') then
			ram(to_integer(unsigned(from_zpu.memAAddr(maxAddrBitBRAM downto 2)))) := from_zpu.memAWrite;
			to_zpu.memARead <= from_zpu.memAWrite;
		else
			to_zpu.memARead <= ram(to_integer(unsigned(from_zpu.memAAddr(maxAddrBitBRAM downto 2))));
		end if;
	end if;
end process;

process (clk)
begin
	if (clk'event and clk = '1') then
		if (from_zpu.memBWriteEnable = '1') then
			ram(to_integer(unsigned(from_zpu.memBAddr(maxAddrBitBRAM downto 2)))) := from_zpu.memBWrite;
			to_zpu.memBRead <= from_zpu.memBWrite;
		else
			to_zpu.memBRead <= ram(to_integer(unsigned(from_zpu.memBAddr(maxAddrBitBRAM downto 2))));
		end if;
	end if;
end process;


end arch;

