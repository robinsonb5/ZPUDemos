-- ZPU
--
-- Copyright 2004-2008 oharboe - �yvind Harboe - oyvind.harboe@zylin.com
-- Modified by Alastair M. Robinson for the ZPUFlex project.
--
-- The FreeBSD license
-- 
-- Redistribution and use in source and binary forms, with or without
-- modification, are permitted provided that the following conditions
-- are met:
-- 
-- 1. Redistributions of source code must retain the above copyright
--    notice, this list of conditions and the following disclaimer.
-- 2. Redistributions in binary form must reproduce the above
--    copyright notice, this list of conditions and the following
--    disclaimer in the documentation and/or other materials
--    provided with the distribution.
-- 
-- THIS SOFTWARE IS PROVIDED BY THE ZPU PROJECT ``AS IS'' AND ANY
-- EXPRESS OR IMPLIED WARRANTIES, INCLUDING, BUT NOT LIMITED TO,
-- THE IMPLIED WARRANTIES OF MERCHANTABILITY AND FITNESS FOR A
-- PARTICULAR PURPOSE ARE DISCLAIMED. IN NO EVENT SHALL THE
-- ZPU PROJECT OR CONTRIBUTORS BE LIABLE FOR ANY DIRECT,
-- INDIRECT, INCIDENTAL, SPECIAL, EXEMPLARY, OR CONSEQUENTIAL DAMAGES
-- (INCLUDING, BUT NOT LIMITED TO, PROCUREMENT OF SUBSTITUTE GOODS
-- OR SERVICES; LOSS OF USE, DATA, OR PROFITS; OR BUSINESS INTERRUPTION)
-- HOWEVER CAUSED AND ON ANY THEORY OF LIABILITY, WHETHER IN CONTRACT,
-- STRICT LIABILITY, OR TORT (INCLUDING NEGLIGENCE OR OTHERWISE)
-- ARISING IN ANY WAY OUT OF THE USE OF THIS SOFTWARE, EVEN IF
-- ADVISED OF THE POSSIBILITY OF SUCH DAMAGE.
-- 
-- The views and conclusions contained in the software and documentation
-- are those of the authors and should not be interpreted as representing
-- official policies, either expressed or implied, of the ZPU Project.

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;


library work;
use work.zpu_config.all;
use work.zpupkg.all;

entity Dhrystone_fast_ROM is
generic
	(
		maxAddrBitBRAM : integer := maxAddrBitBRAMLimit -- Specify your actual ROM size to save LEs and unnecessary block RAM usage.
	);
port (
	clk : in std_logic;
	areset : in std_logic := '0';
	from_zpu : in ZPU_ToROM;
	to_zpu : out ZPU_FromROM
);
end Dhrystone_fast_ROM;

architecture arch of Dhrystone_fast_ROM is

type ram_type is array(natural range 0 to ((2**(maxAddrBitBRAM+1))/4)-1) of std_logic_vector(wordSize-1 downto 0);

shared variable ram : ram_type :=
(
     0 => x"0b0b0b88",
     1 => x"e5040000",
     2 => x"00000000",
     3 => x"00000000",
     4 => x"00000000",
     5 => x"00000000",
     6 => x"00000000",
     7 => x"00000000",
     8 => x"88088c08",
     9 => x"90080b0b",
    10 => x"0b88e108",
    11 => x"2d900c8c",
    12 => x"0c880c04",
    13 => x"00000000",
    14 => x"00000000",
    15 => x"00000000",
    16 => x"71fd0608",
    17 => x"72830609",
    18 => x"81058205",
    19 => x"832b2a83",
    20 => x"ffff0652",
    21 => x"04000000",
    22 => x"00000000",
    23 => x"00000000",
    24 => x"71fd0608",
    25 => x"83ffff73",
    26 => x"83060981",
    27 => x"05820583",
    28 => x"2b2b0906",
    29 => x"7383ffff",
    30 => x"0b0b0b0b",
    31 => x"83a50400",
    32 => x"72098105",
    33 => x"72057373",
    34 => x"09060906",
    35 => x"73097306",
    36 => x"070a8106",
    37 => x"53510400",
    38 => x"00000000",
    39 => x"00000000",
    40 => x"72722473",
    41 => x"732e0753",
    42 => x"51040000",
    43 => x"00000000",
    44 => x"00000000",
    45 => x"00000000",
    46 => x"00000000",
    47 => x"00000000",
    48 => x"71737109",
    49 => x"71068106",
    50 => x"09810572",
    51 => x"0a100a72",
    52 => x"0a100a31",
    53 => x"050a8106",
    54 => x"51515351",
    55 => x"04000000",
    56 => x"72722673",
    57 => x"732e0753",
    58 => x"51040000",
    59 => x"00000000",
    60 => x"00000000",
    61 => x"00000000",
    62 => x"00000000",
    63 => x"00000000",
    64 => x"00000000",
    65 => x"00000000",
    66 => x"00000000",
    67 => x"00000000",
    68 => x"00000000",
    69 => x"00000000",
    70 => x"00000000",
    71 => x"00000000",
    72 => x"0b0b0b88",
    73 => x"ba040000",
    74 => x"00000000",
    75 => x"00000000",
    76 => x"00000000",
    77 => x"00000000",
    78 => x"00000000",
    79 => x"00000000",
    80 => x"720a722b",
    81 => x"0a535104",
    82 => x"00000000",
    83 => x"00000000",
    84 => x"00000000",
    85 => x"00000000",
    86 => x"00000000",
    87 => x"00000000",
    88 => x"72729f06",
    89 => x"0981050b",
    90 => x"0b0b889f",
    91 => x"05040000",
    92 => x"00000000",
    93 => x"00000000",
    94 => x"00000000",
    95 => x"00000000",
    96 => x"72722aff",
    97 => x"739f062a",
    98 => x"0974090a",
    99 => x"8106ff05",
   100 => x"06075351",
   101 => x"04000000",
   102 => x"00000000",
   103 => x"00000000",
   104 => x"71715351",
   105 => x"04067383",
   106 => x"06098105",
   107 => x"8205832b",
   108 => x"0b2b0772",
   109 => x"fc060c51",
   110 => x"51040000",
   111 => x"00000000",
   112 => x"72098105",
   113 => x"72050970",
   114 => x"81050906",
   115 => x"0a810653",
   116 => x"51040000",
   117 => x"00000000",
   118 => x"00000000",
   119 => x"00000000",
   120 => x"72098105",
   121 => x"72050970",
   122 => x"81050906",
   123 => x"0a098106",
   124 => x"53510400",
   125 => x"00000000",
   126 => x"00000000",
   127 => x"00000000",
   128 => x"71098105",
   129 => x"52040000",
   130 => x"00000000",
   131 => x"00000000",
   132 => x"00000000",
   133 => x"00000000",
   134 => x"00000000",
   135 => x"00000000",
   136 => x"72720981",
   137 => x"05055351",
   138 => x"04000000",
   139 => x"00000000",
   140 => x"00000000",
   141 => x"00000000",
   142 => x"00000000",
   143 => x"00000000",
   144 => x"72097206",
   145 => x"73730906",
   146 => x"07535104",
   147 => x"00000000",
   148 => x"00000000",
   149 => x"00000000",
   150 => x"00000000",
   151 => x"00000000",
   152 => x"71fc0608",
   153 => x"72830609",
   154 => x"81058305",
   155 => x"1010102a",
   156 => x"81ff0652",
   157 => x"04000000",
   158 => x"00000000",
   159 => x"00000000",
   160 => x"71fc0608",
   161 => x"0b0b0ba2",
   162 => x"b4738306",
   163 => x"10100508",
   164 => x"060b0b0b",
   165 => x"88a20400",
   166 => x"00000000",
   167 => x"00000000",
   168 => x"88088c08",
   169 => x"90087575",
   170 => x"0b0b0b9b",
   171 => x"a82d5050",
   172 => x"88085690",
   173 => x"0c8c0c88",
   174 => x"0c510400",
   175 => x"00000000",
   176 => x"88088c08",
   177 => x"90087575",
   178 => x"0b0b0b9c",
   179 => x"da2d5050",
   180 => x"88085690",
   181 => x"0c8c0c88",
   182 => x"0c510400",
   183 => x"00000000",
   184 => x"72097081",
   185 => x"0509060a",
   186 => x"8106ff05",
   187 => x"70547106",
   188 => x"73097274",
   189 => x"05ff0506",
   190 => x"07515151",
   191 => x"04000000",
   192 => x"72097081",
   193 => x"0509060a",
   194 => x"098106ff",
   195 => x"05705471",
   196 => x"06730972",
   197 => x"7405ff05",
   198 => x"06075151",
   199 => x"51040000",
   200 => x"05ff0504",
   201 => x"00000000",
   202 => x"00000000",
   203 => x"00000000",
   204 => x"00000000",
   205 => x"00000000",
   206 => x"00000000",
   207 => x"00000000",
   208 => x"04000000",
   209 => x"00000000",
   210 => x"00000000",
   211 => x"00000000",
   212 => x"00000000",
   213 => x"00000000",
   214 => x"00000000",
   215 => x"00000000",
   216 => x"71810552",
   217 => x"04000000",
   218 => x"00000000",
   219 => x"00000000",
   220 => x"00000000",
   221 => x"00000000",
   222 => x"00000000",
   223 => x"00000000",
   224 => x"00000000",
   225 => x"00000000",
   226 => x"00000000",
   227 => x"00000000",
   228 => x"00000000",
   229 => x"00000000",
   230 => x"00000000",
   231 => x"00000000",
   232 => x"02840572",
   233 => x"10100552",
   234 => x"04000000",
   235 => x"00000000",
   236 => x"00000000",
   237 => x"00000000",
   238 => x"00000000",
   239 => x"00000000",
   240 => x"00000000",
   241 => x"00000000",
   242 => x"00000000",
   243 => x"00000000",
   244 => x"00000000",
   245 => x"00000000",
   246 => x"00000000",
   247 => x"00000000",
   248 => x"717105ff",
   249 => x"05715351",
   250 => x"020d0400",
   251 => x"00000000",
   252 => x"00000000",
   253 => x"00000000",
   254 => x"00000000",
   255 => x"00000000",
   256 => x"10101010",
   257 => x"10101010",
   258 => x"10101010",
   259 => x"10101010",
   260 => x"10101010",
   261 => x"10101010",
   262 => x"10101010",
   263 => x"10101053",
   264 => x"51047381",
   265 => x"ff067383",
   266 => x"06098105",
   267 => x"83051010",
   268 => x"102b0772",
   269 => x"fc060c51",
   270 => x"51047272",
   271 => x"80728106",
   272 => x"ff050972",
   273 => x"06057110",
   274 => x"52720a10",
   275 => x"0a5372ed",
   276 => x"38515153",
   277 => x"51040000",
   278 => x"800488da",
   279 => x"04040000",
   280 => x"00000004",
   281 => x"5d88da0b",
   282 => x"91a00402",
   283 => x"c0050d02",
   284 => x"80c4055b",
   285 => x"80707c70",
   286 => x"84055e08",
   287 => x"725f5f5f",
   288 => x"587c7084",
   289 => x"055e0857",
   290 => x"80597698",
   291 => x"2a77882b",
   292 => x"58557480",
   293 => x"2e848d38",
   294 => x"7b802e80",
   295 => x"c838805c",
   296 => x"7480e42e",
   297 => x"81f93874",
   298 => x"80f82e81",
   299 => x"f2387480",
   300 => x"e42e81fd",
   301 => x"387480e4",
   302 => x"2680dd38",
   303 => x"7480e32e",
   304 => x"bb38a551",
   305 => x"8ddd2d74",
   306 => x"518ddd2d",
   307 => x"82185881",
   308 => x"19598379",
   309 => x"25ffb338",
   310 => x"74ffa638",
   311 => x"7e880c02",
   312 => x"80c0050d",
   313 => x"0474a52e",
   314 => x"09810698",
   315 => x"38810b81",
   316 => x"1a5a5c83",
   317 => x"7925ff92",
   318 => x"3889d804",
   319 => x"7a841c71",
   320 => x"08575c56",
   321 => x"74518ddd",
   322 => x"2d811881",
   323 => x"1a5a5883",
   324 => x"7925fef6",
   325 => x"3889d804",
   326 => x"7480f32e",
   327 => x"838f3874",
   328 => x"80f82e09",
   329 => x"8106ff9a",
   330 => x"387d0b0b",
   331 => x"0ba7dc0b",
   332 => x"0b0b0ba7",
   333 => x"8c565b53",
   334 => x"8056757e",
   335 => x"24839138",
   336 => x"7281c538",
   337 => x"b00b0b0b",
   338 => x"0ba78c0b",
   339 => x"85802d81",
   340 => x"1454ff14",
   341 => x"547384e0",
   342 => x"2d7a7081",
   343 => x"055c8580",
   344 => x"2d811656",
   345 => x"730b0b0b",
   346 => x"a78c2e09",
   347 => x"8106e338",
   348 => x"807a8580",
   349 => x"2d750b0b",
   350 => x"0ba7dc57",
   351 => x"53ff1354",
   352 => x"807325fe",
   353 => x"ca387570",
   354 => x"81055784",
   355 => x"e02d7052",
   356 => x"558ddd2d",
   357 => x"811874ff",
   358 => x"16565458",
   359 => x"8b80047a",
   360 => x"841c7108",
   361 => x"405c5374",
   362 => x"80e42e09",
   363 => x"8106fe85",
   364 => x"387d0b0b",
   365 => x"0ba7dc0b",
   366 => x"0b0b0ba7",
   367 => x"8c565b53",
   368 => x"8056757e",
   369 => x"2481fc38",
   370 => x"72818b38",
   371 => x"b00b0b0b",
   372 => x"0ba78c0b",
   373 => x"85802d81",
   374 => x"1454ff14",
   375 => x"547384e0",
   376 => x"2d7a7081",
   377 => x"055c8580",
   378 => x"2d811656",
   379 => x"730b0b0b",
   380 => x"a78c2e09",
   381 => x"8106e338",
   382 => x"807a8580",
   383 => x"2d750b0b",
   384 => x"0ba7dc57",
   385 => x"538afd04",
   386 => x"90527251",
   387 => x"9cda2d88",
   388 => x"08a2c405",
   389 => x"84e02d74",
   390 => x"70810556",
   391 => x"85802d90",
   392 => x"5272519b",
   393 => x"a82d8808",
   394 => x"538808dc",
   395 => x"38730b0b",
   396 => x"0ba78c2e",
   397 => x"feba38ff",
   398 => x"14547384",
   399 => x"e02d7a70",
   400 => x"81055c85",
   401 => x"802d8116",
   402 => x"56730b0b",
   403 => x"0ba78c2e",
   404 => x"fe9e388a",
   405 => x"d2048a52",
   406 => x"72519cda",
   407 => x"2d8808a2",
   408 => x"c40584e0",
   409 => x"2d747081",
   410 => x"05568580",
   411 => x"2d8a5272",
   412 => x"519ba82d",
   413 => x"88085388",
   414 => x"08dc3873",
   415 => x"0b0b0ba7",
   416 => x"8c2efdec",
   417 => x"38ff1454",
   418 => x"7384e02d",
   419 => x"7a708105",
   420 => x"5c85802d",
   421 => x"81165673",
   422 => x"0b0b0ba7",
   423 => x"8c2efed8",
   424 => x"388bda04",
   425 => x"77880c02",
   426 => x"80c0050d",
   427 => x"047a841c",
   428 => x"71087054",
   429 => x"585c548d",
   430 => x"fe2d800b",
   431 => x"ff115553",
   432 => x"8b8004ad",
   433 => x"518ddd2d",
   434 => x"7d098105",
   435 => x"538bc804",
   436 => x"ad518ddd",
   437 => x"2d7d0981",
   438 => x"05538ac0",
   439 => x"0402f805",
   440 => x"0d7352c0",
   441 => x"0870882a",
   442 => x"70810651",
   443 => x"51517080",
   444 => x"2ef13871",
   445 => x"c00c7188",
   446 => x"0c028805",
   447 => x"0d0402e8",
   448 => x"050d8078",
   449 => x"57557570",
   450 => x"84055708",
   451 => x"53805472",
   452 => x"982a7388",
   453 => x"2b545271",
   454 => x"802ea238",
   455 => x"c0087088",
   456 => x"2a708106",
   457 => x"51515170",
   458 => x"802ef138",
   459 => x"71c00c81",
   460 => x"15811555",
   461 => x"55837425",
   462 => x"d63871ca",
   463 => x"3874880c",
   464 => x"0298050d",
   465 => x"04c80888",
   466 => x"0c0402fc",
   467 => x"050d80c1",
   468 => x"0b80f7a8",
   469 => x"0b85802d",
   470 => x"800b80f9",
   471 => x"c00c7088",
   472 => x"0c028405",
   473 => x"0d0402f8",
   474 => x"050d800b",
   475 => x"80f7a80b",
   476 => x"84e02d52",
   477 => x"527080c1",
   478 => x"2e9d3871",
   479 => x"80f9c008",
   480 => x"0780f9c0",
   481 => x"0c80c20b",
   482 => x"80f7ac0b",
   483 => x"85802d70",
   484 => x"880c0288",
   485 => x"050d0481",
   486 => x"0b80f9c0",
   487 => x"080780f9",
   488 => x"c00c80c2",
   489 => x"0b80f7ac",
   490 => x"0b85802d",
   491 => x"70880c02",
   492 => x"88050d04",
   493 => x"02f0050d",
   494 => x"7570088a",
   495 => x"05535380",
   496 => x"f7a80b84",
   497 => x"e02d5170",
   498 => x"80c12e8c",
   499 => x"3873f038",
   500 => x"70880c02",
   501 => x"90050d04",
   502 => x"ff127080",
   503 => x"f7a40831",
   504 => x"740c880c",
   505 => x"0290050d",
   506 => x"0402ec05",
   507 => x"0d80f7d0",
   508 => x"08557480",
   509 => x"2e8c3876",
   510 => x"7508710c",
   511 => x"80f7d008",
   512 => x"56548c15",
   513 => x"5380f7a4",
   514 => x"08528a51",
   515 => x"98fe2d73",
   516 => x"880c0294",
   517 => x"050d0402",
   518 => x"e8050d77",
   519 => x"70085656",
   520 => x"b05380f7",
   521 => x"d0085274",
   522 => x"51a0862d",
   523 => x"850b8c17",
   524 => x"0c850b8c",
   525 => x"160c7508",
   526 => x"750c80f7",
   527 => x"d0085473",
   528 => x"802e8a38",
   529 => x"7308750c",
   530 => x"80f7d008",
   531 => x"548c1453",
   532 => x"80f7a408",
   533 => x"528a5198",
   534 => x"fe2d8415",
   535 => x"08ae3886",
   536 => x"0b8c160c",
   537 => x"88155288",
   538 => x"16085198",
   539 => x"982d80f7",
   540 => x"d0087008",
   541 => x"760c548c",
   542 => x"15705454",
   543 => x"8a527308",
   544 => x"5198fe2d",
   545 => x"73880c02",
   546 => x"98050d04",
   547 => x"750854b0",
   548 => x"53735275",
   549 => x"51a0862d",
   550 => x"73880c02",
   551 => x"98050d04",
   552 => x"02c8050d",
   553 => x"80f6bc0b",
   554 => x"80f6f00c",
   555 => x"80f6f40b",
   556 => x"80f7d00c",
   557 => x"80f6bc0b",
   558 => x"80f6f40c",
   559 => x"800b80f6",
   560 => x"f40b8405",
   561 => x"0c820b80",
   562 => x"f6f40b88",
   563 => x"050ca80b",
   564 => x"80f6f40b",
   565 => x"8c050c9f",
   566 => x"53a2d852",
   567 => x"80f78451",
   568 => x"a0862d9f",
   569 => x"53a2f852",
   570 => x"80f9a051",
   571 => x"a0862d8a",
   572 => x"0bb5880c",
   573 => x"a5d85188",
   574 => x"eb2da398",
   575 => x"5188eb2d",
   576 => x"a5d85188",
   577 => x"eb2da788",
   578 => x"08802e84",
   579 => x"9138a3c8",
   580 => x"5188eb2d",
   581 => x"a5d85188",
   582 => x"eb2da784",
   583 => x"0852a3f4",
   584 => x"5188eb2d",
   585 => x"c80870a8",
   586 => x"a80c5681",
   587 => x"58800ba7",
   588 => x"84082582",
   589 => x"dc3802ac",
   590 => x"055b80c1",
   591 => x"0b80f7a8",
   592 => x"0b85802d",
   593 => x"810b80f9",
   594 => x"c00c80c2",
   595 => x"0b80f7ac",
   596 => x"0b85802d",
   597 => x"825c835a",
   598 => x"9f53a4a4",
   599 => x"5280f7b0",
   600 => x"51a0862d",
   601 => x"815d800b",
   602 => x"80f7b053",
   603 => x"80f9a052",
   604 => x"559ab02d",
   605 => x"8808752e",
   606 => x"09810683",
   607 => x"38815574",
   608 => x"80f9c00c",
   609 => x"7b705755",
   610 => x"748325a1",
   611 => x"38741010",
   612 => x"15fd055e",
   613 => x"02b805fc",
   614 => x"05538352",
   615 => x"755198fe",
   616 => x"2d811c70",
   617 => x"5d705755",
   618 => x"837524e1",
   619 => x"387d5474",
   620 => x"53a8ac52",
   621 => x"80f7d851",
   622 => x"99902d80",
   623 => x"f7d00870",
   624 => x"085757b0",
   625 => x"53765275",
   626 => x"51a0862d",
   627 => x"850b8c18",
   628 => x"0c850b8c",
   629 => x"170c7608",
   630 => x"760c80f7",
   631 => x"d0085574",
   632 => x"802e8a38",
   633 => x"7408760c",
   634 => x"80f7d008",
   635 => x"558c1553",
   636 => x"80f7a408",
   637 => x"528a5198",
   638 => x"fe2d8416",
   639 => x"0883d838",
   640 => x"860b8c17",
   641 => x"0c881652",
   642 => x"88170851",
   643 => x"98982d80",
   644 => x"f7d00870",
   645 => x"08770c57",
   646 => x"8c167054",
   647 => x"558a5274",
   648 => x"085198fe",
   649 => x"2d80c10b",
   650 => x"80f7ac0b",
   651 => x"84e02d56",
   652 => x"56757526",
   653 => x"a53880c3",
   654 => x"52755199",
   655 => x"fc2d8808",
   656 => x"7d2e82e2",
   657 => x"38811670",
   658 => x"81ff0680",
   659 => x"f7ac0b84",
   660 => x"e02d5257",
   661 => x"55747627",
   662 => x"dd38797c",
   663 => x"297e5351",
   664 => x"9ba82d88",
   665 => x"085c8808",
   666 => x"8a0580f7",
   667 => x"a80b84e0",
   668 => x"2d80f7a4",
   669 => x"08595755",
   670 => x"7580c12e",
   671 => x"82f43878",
   672 => x"f7388118",
   673 => x"58a78408",
   674 => x"7825fdae",
   675 => x"38a8a808",
   676 => x"56c80870",
   677 => x"80f6ec0c",
   678 => x"70773170",
   679 => x"a8a40c53",
   680 => x"a4c4525b",
   681 => x"88eb2da8",
   682 => x"a4085680",
   683 => x"f7762580",
   684 => x"f338a784",
   685 => x"08705376",
   686 => x"87e82952",
   687 => x"5a9ba82d",
   688 => x"8808a89c",
   689 => x"0c755279",
   690 => x"87e82951",
   691 => x"9ba82d88",
   692 => x"08a8a00c",
   693 => x"75527984",
   694 => x"b929519b",
   695 => x"a82d8808",
   696 => x"80f7d40c",
   697 => x"a4d45188",
   698 => x"eb2da89c",
   699 => x"0852a584",
   700 => x"5188eb2d",
   701 => x"a58c5188",
   702 => x"eb2da8a0",
   703 => x"0852a584",
   704 => x"5188eb2d",
   705 => x"80f7d408",
   706 => x"52a5bc51",
   707 => x"88eb2da5",
   708 => x"d85188eb",
   709 => x"2d800b88",
   710 => x"0c02b805",
   711 => x"0d04a5dc",
   712 => x"51929104",
   713 => x"a68c5188",
   714 => x"eb2da6c4",
   715 => x"5188eb2d",
   716 => x"a5d85188",
   717 => x"eb2da8a4",
   718 => x"08a78408",
   719 => x"70547187",
   720 => x"e829535b",
   721 => x"569ba82d",
   722 => x"8808a89c",
   723 => x"0c755279",
   724 => x"87e82951",
   725 => x"9ba82d88",
   726 => x"08a8a00c",
   727 => x"75527984",
   728 => x"b929519b",
   729 => x"a82d8808",
   730 => x"80f7d40c",
   731 => x"a4d45188",
   732 => x"eb2da89c",
   733 => x"0852a584",
   734 => x"5188eb2d",
   735 => x"a58c5188",
   736 => x"eb2da8a0",
   737 => x"0852a584",
   738 => x"5188eb2d",
   739 => x"80f7d408",
   740 => x"52a5bc51",
   741 => x"88eb2da5",
   742 => x"d85188eb",
   743 => x"2d800b88",
   744 => x"0c02b805",
   745 => x"0d0402b8",
   746 => x"05f80552",
   747 => x"80519898",
   748 => x"2d9f53a6",
   749 => x"e45280f7",
   750 => x"b051a086",
   751 => x"2d777880",
   752 => x"f7a40c81",
   753 => x"177081ff",
   754 => x"0680f7ac",
   755 => x"0b84e02d",
   756 => x"5258565a",
   757 => x"94d50476",
   758 => x"0856b053",
   759 => x"75527651",
   760 => x"a0862d80",
   761 => x"c10b80f7",
   762 => x"ac0b84e0",
   763 => x"2d565694",
   764 => x"b104ff15",
   765 => x"7078317c",
   766 => x"0c598059",
   767 => x"95820402",
   768 => x"f8050d73",
   769 => x"82327009",
   770 => x"81057072",
   771 => x"07802588",
   772 => x"0c525202",
   773 => x"88050d04",
   774 => x"02f4050d",
   775 => x"74767153",
   776 => x"54527182",
   777 => x"2e833883",
   778 => x"5171812e",
   779 => x"9b388172",
   780 => x"26a03871",
   781 => x"822ebc38",
   782 => x"71842eac",
   783 => x"3870730c",
   784 => x"70880c02",
   785 => x"8c050d04",
   786 => x"80e40b80",
   787 => x"f7a40825",
   788 => x"8c388073",
   789 => x"0c70880c",
   790 => x"028c050d",
   791 => x"0483730c",
   792 => x"70880c02",
   793 => x"8c050d04",
   794 => x"82730c70",
   795 => x"880c028c",
   796 => x"050d0481",
   797 => x"730c7088",
   798 => x"0c028c05",
   799 => x"0d0402fc",
   800 => x"050d7474",
   801 => x"14820571",
   802 => x"0c880c02",
   803 => x"84050d04",
   804 => x"02d8050d",
   805 => x"7b7d7f61",
   806 => x"85127082",
   807 => x"2b751170",
   808 => x"74717084",
   809 => x"05530c5a",
   810 => x"5a5d5b76",
   811 => x"0c7980f8",
   812 => x"180c7986",
   813 => x"12525758",
   814 => x"5a5a7676",
   815 => x"24993876",
   816 => x"b329822b",
   817 => x"79115153",
   818 => x"76737084",
   819 => x"05550c81",
   820 => x"14547574",
   821 => x"25f23876",
   822 => x"81cc2919",
   823 => x"fc110881",
   824 => x"05fc120c",
   825 => x"7a197008",
   826 => x"9fa0130c",
   827 => x"5856850b",
   828 => x"80f7a40c",
   829 => x"75880c02",
   830 => x"a8050d04",
   831 => x"02f4050d",
   832 => x"02930584",
   833 => x"e02d5180",
   834 => x"02840597",
   835 => x"0584e02d",
   836 => x"54527073",
   837 => x"2e893871",
   838 => x"880c028c",
   839 => x"050d0470",
   840 => x"80f7a80b",
   841 => x"85802d81",
   842 => x"0b880c02",
   843 => x"8c050d04",
   844 => x"02dc050d",
   845 => x"7a7c5956",
   846 => x"820b8319",
   847 => x"55557416",
   848 => x"7084e02d",
   849 => x"7584e02d",
   850 => x"5b515372",
   851 => x"792e80c7",
   852 => x"3880c10b",
   853 => x"81168116",
   854 => x"56565782",
   855 => x"7525df38",
   856 => x"ffa91770",
   857 => x"81ff0655",
   858 => x"59738226",
   859 => x"83388755",
   860 => x"81537680",
   861 => x"d22e9838",
   862 => x"77527551",
   863 => x"a19f2d80",
   864 => x"53728808",
   865 => x"25893887",
   866 => x"1580f7a4",
   867 => x"0c815372",
   868 => x"880c02a4",
   869 => x"050d0472",
   870 => x"80f7a80b",
   871 => x"85802d82",
   872 => x"7525ff9a",
   873 => x"389ae004",
   874 => x"94080294",
   875 => x"0cf93d0d",
   876 => x"800b9408",
   877 => x"fc050c94",
   878 => x"08880508",
   879 => x"8025ab38",
   880 => x"94088805",
   881 => x"08309408",
   882 => x"88050c80",
   883 => x"0b9408f4",
   884 => x"050c9408",
   885 => x"fc050888",
   886 => x"38810b94",
   887 => x"08f4050c",
   888 => x"9408f405",
   889 => x"089408fc",
   890 => x"050c9408",
   891 => x"8c050880",
   892 => x"25ab3894",
   893 => x"088c0508",
   894 => x"3094088c",
   895 => x"050c800b",
   896 => x"9408f005",
   897 => x"0c9408fc",
   898 => x"05088838",
   899 => x"810b9408",
   900 => x"f0050c94",
   901 => x"08f00508",
   902 => x"9408fc05",
   903 => x"0c805394",
   904 => x"088c0508",
   905 => x"52940888",
   906 => x"05085181",
   907 => x"a73f8808",
   908 => x"709408f8",
   909 => x"050c5494",
   910 => x"08fc0508",
   911 => x"802e8c38",
   912 => x"9408f805",
   913 => x"08309408",
   914 => x"f8050c94",
   915 => x"08f80508",
   916 => x"70880c54",
   917 => x"893d0d94",
   918 => x"0c049408",
   919 => x"02940cfb",
   920 => x"3d0d800b",
   921 => x"9408fc05",
   922 => x"0c940888",
   923 => x"05088025",
   924 => x"93389408",
   925 => x"88050830",
   926 => x"94088805",
   927 => x"0c810b94",
   928 => x"08fc050c",
   929 => x"94088c05",
   930 => x"0880258c",
   931 => x"3894088c",
   932 => x"05083094",
   933 => x"088c050c",
   934 => x"81539408",
   935 => x"8c050852",
   936 => x"94088805",
   937 => x"0851ad3f",
   938 => x"88087094",
   939 => x"08f8050c",
   940 => x"549408fc",
   941 => x"0508802e",
   942 => x"8c389408",
   943 => x"f8050830",
   944 => x"9408f805",
   945 => x"0c9408f8",
   946 => x"05087088",
   947 => x"0c54873d",
   948 => x"0d940c04",
   949 => x"94080294",
   950 => x"0cfd3d0d",
   951 => x"810b9408",
   952 => x"fc050c80",
   953 => x"0b9408f8",
   954 => x"050c9408",
   955 => x"8c050894",
   956 => x"08880508",
   957 => x"27ac3894",
   958 => x"08fc0508",
   959 => x"802ea338",
   960 => x"800b9408",
   961 => x"8c050824",
   962 => x"99389408",
   963 => x"8c050810",
   964 => x"94088c05",
   965 => x"0c9408fc",
   966 => x"05081094",
   967 => x"08fc050c",
   968 => x"c9399408",
   969 => x"fc050880",
   970 => x"2e80c938",
   971 => x"94088c05",
   972 => x"08940888",
   973 => x"050826a1",
   974 => x"38940888",
   975 => x"05089408",
   976 => x"8c050831",
   977 => x"94088805",
   978 => x"0c9408f8",
   979 => x"05089408",
   980 => x"fc050807",
   981 => x"9408f805",
   982 => x"0c9408fc",
   983 => x"0508812a",
   984 => x"9408fc05",
   985 => x"0c94088c",
   986 => x"0508812a",
   987 => x"94088c05",
   988 => x"0cffaf39",
   989 => x"94089005",
   990 => x"08802e8f",
   991 => x"38940888",
   992 => x"05087094",
   993 => x"08f4050c",
   994 => x"518d3994",
   995 => x"08f80508",
   996 => x"709408f4",
   997 => x"050c5194",
   998 => x"08f40508",
   999 => x"880c853d",
  1000 => x"0d940c04",
  1001 => x"94080294",
  1002 => x"0cff3d0d",
  1003 => x"800b9408",
  1004 => x"fc050c94",
  1005 => x"08880508",
  1006 => x"8106ff11",
  1007 => x"70097094",
  1008 => x"088c0508",
  1009 => x"069408fc",
  1010 => x"05081194",
  1011 => x"08fc050c",
  1012 => x"94088805",
  1013 => x"08812a94",
  1014 => x"0888050c",
  1015 => x"94088c05",
  1016 => x"08109408",
  1017 => x"8c050c51",
  1018 => x"51515194",
  1019 => x"08880508",
  1020 => x"802e8438",
  1021 => x"ffbd3994",
  1022 => x"08fc0508",
  1023 => x"70880c51",
  1024 => x"833d0d94",
  1025 => x"0c04fc3d",
  1026 => x"0d767079",
  1027 => x"7b555555",
  1028 => x"558f7227",
  1029 => x"8c387275",
  1030 => x"07830651",
  1031 => x"70802ea7",
  1032 => x"38ff1252",
  1033 => x"71ff2e98",
  1034 => x"38727081",
  1035 => x"05543374",
  1036 => x"70810556",
  1037 => x"34ff1252",
  1038 => x"71ff2e09",
  1039 => x"8106ea38",
  1040 => x"74880c86",
  1041 => x"3d0d0474",
  1042 => x"51727084",
  1043 => x"05540871",
  1044 => x"70840553",
  1045 => x"0c727084",
  1046 => x"05540871",
  1047 => x"70840553",
  1048 => x"0c727084",
  1049 => x"05540871",
  1050 => x"70840553",
  1051 => x"0c727084",
  1052 => x"05540871",
  1053 => x"70840553",
  1054 => x"0cf01252",
  1055 => x"718f26c9",
  1056 => x"38837227",
  1057 => x"95387270",
  1058 => x"84055408",
  1059 => x"71708405",
  1060 => x"530cfc12",
  1061 => x"52718326",
  1062 => x"ed387054",
  1063 => x"ff8339fb",
  1064 => x"3d0d7779",
  1065 => x"70720783",
  1066 => x"06535452",
  1067 => x"70933871",
  1068 => x"73730854",
  1069 => x"56547173",
  1070 => x"082e80c4",
  1071 => x"38737554",
  1072 => x"52713370",
  1073 => x"81ff0652",
  1074 => x"5470802e",
  1075 => x"9d387233",
  1076 => x"5570752e",
  1077 => x"09810695",
  1078 => x"38811281",
  1079 => x"14713370",
  1080 => x"81ff0654",
  1081 => x"56545270",
  1082 => x"e5387233",
  1083 => x"557381ff",
  1084 => x"067581ff",
  1085 => x"06717131",
  1086 => x"880c5252",
  1087 => x"873d0d04",
  1088 => x"710970f7",
  1089 => x"fbfdff14",
  1090 => x"0670f884",
  1091 => x"82818006",
  1092 => x"51515170",
  1093 => x"97388414",
  1094 => x"84167108",
  1095 => x"54565471",
  1096 => x"75082edc",
  1097 => x"38737554",
  1098 => x"52ff9639",
  1099 => x"800b880c",
  1100 => x"873d0d04",
  1101 => x"00ffffff",
  1102 => x"ff00ffff",
  1103 => x"ffff00ff",
  1104 => x"ffffff00",
  1105 => x"30313233",
  1106 => x"34353637",
  1107 => x"38394142",
  1108 => x"43444546",
  1109 => x"00000000",
  1110 => x"44485259",
  1111 => x"53544f4e",
  1112 => x"45205052",
  1113 => x"4f475241",
  1114 => x"4d2c2053",
  1115 => x"4f4d4520",
  1116 => x"53545249",
  1117 => x"4e470000",
  1118 => x"44485259",
  1119 => x"53544f4e",
  1120 => x"45205052",
  1121 => x"4f475241",
  1122 => x"4d2c2031",
  1123 => x"27535420",
  1124 => x"53545249",
  1125 => x"4e470000",
  1126 => x"44687279",
  1127 => x"73746f6e",
  1128 => x"65204265",
  1129 => x"6e63686d",
  1130 => x"61726b2c",
  1131 => x"20566572",
  1132 => x"73696f6e",
  1133 => x"20322e31",
  1134 => x"20284c61",
  1135 => x"6e677561",
  1136 => x"67653a20",
  1137 => x"43290a00",
  1138 => x"50726f67",
  1139 => x"72616d20",
  1140 => x"636f6d70",
  1141 => x"696c6564",
  1142 => x"20776974",
  1143 => x"68202772",
  1144 => x"65676973",
  1145 => x"74657227",
  1146 => x"20617474",
  1147 => x"72696275",
  1148 => x"74650a00",
  1149 => x"45786563",
  1150 => x"7574696f",
  1151 => x"6e207374",
  1152 => x"61727473",
  1153 => x"2c202564",
  1154 => x"2072756e",
  1155 => x"73207468",
  1156 => x"726f7567",
  1157 => x"68204468",
  1158 => x"72797374",
  1159 => x"6f6e650a",
  1160 => x"00000000",
  1161 => x"44485259",
  1162 => x"53544f4e",
  1163 => x"45205052",
  1164 => x"4f475241",
  1165 => x"4d2c2032",
  1166 => x"274e4420",
  1167 => x"53545249",
  1168 => x"4e470000",
  1169 => x"55736572",
  1170 => x"2074696d",
  1171 => x"653a2025",
  1172 => x"640a0000",
  1173 => x"4d696372",
  1174 => x"6f736563",
  1175 => x"6f6e6473",
  1176 => x"20666f72",
  1177 => x"206f6e65",
  1178 => x"2072756e",
  1179 => x"20746872",
  1180 => x"6f756768",
  1181 => x"20446872",
  1182 => x"7973746f",
  1183 => x"6e653a20",
  1184 => x"00000000",
  1185 => x"2564200a",
  1186 => x"00000000",
  1187 => x"44687279",
  1188 => x"73746f6e",
  1189 => x"65732070",
  1190 => x"65722053",
  1191 => x"65636f6e",
  1192 => x"643a2020",
  1193 => x"20202020",
  1194 => x"20202020",
  1195 => x"20202020",
  1196 => x"20202020",
  1197 => x"20202020",
  1198 => x"00000000",
  1199 => x"56415820",
  1200 => x"4d495053",
  1201 => x"20726174",
  1202 => x"696e6720",
  1203 => x"2a203130",
  1204 => x"3030203d",
  1205 => x"20256420",
  1206 => x"0a000000",
  1207 => x"50726f67",
  1208 => x"72616d20",
  1209 => x"636f6d70",
  1210 => x"696c6564",
  1211 => x"20776974",
  1212 => x"686f7574",
  1213 => x"20277265",
  1214 => x"67697374",
  1215 => x"65722720",
  1216 => x"61747472",
  1217 => x"69627574",
  1218 => x"650a0000",
  1219 => x"4d656173",
  1220 => x"75726564",
  1221 => x"2074696d",
  1222 => x"6520746f",
  1223 => x"6f20736d",
  1224 => x"616c6c20",
  1225 => x"746f206f",
  1226 => x"62746169",
  1227 => x"6e206d65",
  1228 => x"616e696e",
  1229 => x"6766756c",
  1230 => x"20726573",
  1231 => x"756c7473",
  1232 => x"0a000000",
  1233 => x"506c6561",
  1234 => x"73652069",
  1235 => x"6e637265",
  1236 => x"61736520",
  1237 => x"6e756d62",
  1238 => x"6572206f",
  1239 => x"66207275",
  1240 => x"6e730a00",
  1241 => x"44485259",
  1242 => x"53544f4e",
  1243 => x"45205052",
  1244 => x"4f475241",
  1245 => x"4d2c2033",
  1246 => x"27524420",
  1247 => x"53545249",
  1248 => x"4e470000",
  1249 => x"000061a8",
  1250 => x"00000000",
	others => x"00000000"
);

begin

process (clk)
begin
	if (clk'event and clk = '1') then
		if (from_zpu.memAWriteEnable = '1') and (from_zpu.memBWriteEnable = '1') and (from_zpu.memAAddr=from_zpu.memBAddr) and (from_zpu.memAWrite/=from_zpu.memBWrite) then
			report "write collision" severity failure;
		end if;
	
		if (from_zpu.memAWriteEnable = '1') then
			ram(to_integer(unsigned(from_zpu.memAAddr(maxAddrBitBRAM downto 2)))) := from_zpu.memAWrite;
			to_zpu.memARead <= from_zpu.memAWrite;
		else
			to_zpu.memARead <= ram(to_integer(unsigned(from_zpu.memAAddr(maxAddrBitBRAM downto 2))));
		end if;
	end if;
end process;

process (clk)
begin
	if (clk'event and clk = '1') then
		if (from_zpu.memBWriteEnable = '1') then
			ram(to_integer(unsigned(from_zpu.memBAddr(maxAddrBitBRAM downto 2)))) := from_zpu.memBWrite;
			to_zpu.memBRead <= from_zpu.memBWrite;
		else
			to_zpu.memBRead <= ram(to_integer(unsigned(from_zpu.memBAddr(maxAddrBitBRAM downto 2))));
		end if;
	end if;
end process;


end arch;

