-- ZPU
--
-- Copyright 2004-2008 oharboe - �yvind Harboe - oyvind.harboe@zylin.com
-- Modified by Alastair M. Robinson for the ZPUFlex project.
--
-- The FreeBSD license
-- 
-- Redistribution and use in source and binary forms, with or without
-- modification, are permitted provided that the following conditions
-- are met:
-- 
-- 1. Redistributions of source code must retain the above copyright
--    notice, this list of conditions and the following disclaimer.
-- 2. Redistributions in binary form must reproduce the above
--    copyright notice, this list of conditions and the following
--    disclaimer in the documentation and/or other materials
--    provided with the distribution.
-- 
-- THIS SOFTWARE IS PROVIDED BY THE ZPU PROJECT ``AS IS'' AND ANY
-- EXPRESS OR IMPLIED WARRANTIES, INCLUDING, BUT NOT LIMITED TO,
-- THE IMPLIED WARRANTIES OF MERCHANTABILITY AND FITNESS FOR A
-- PARTICULAR PURPOSE ARE DISCLAIMED. IN NO EVENT SHALL THE
-- ZPU PROJECT OR CONTRIBUTORS BE LIABLE FOR ANY DIRECT,
-- INDIRECT, INCIDENTAL, SPECIAL, EXEMPLARY, OR CONSEQUENTIAL DAMAGES
-- (INCLUDING, BUT NOT LIMITED TO, PROCUREMENT OF SUBSTITUTE GOODS
-- OR SERVICES; LOSS OF USE, DATA, OR PROFITS; OR BUSINESS INTERRUPTION)
-- HOWEVER CAUSED AND ON ANY THEORY OF LIABILITY, WHETHER IN CONTRACT,
-- STRICT LIABILITY, OR TORT (INCLUDING NEGLIGENCE OR OTHERWISE)
-- ARISING IN ANY WAY OUT OF THE USE OF THIS SOFTWARE, EVEN IF
-- ADVISED OF THE POSSIBILITY OF SUCH DAMAGE.
-- 
-- The views and conclusions contained in the software and documentation
-- are those of the authors and should not be interpreted as representing
-- official policies, either expressed or implied, of the ZPU Project.

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;


library work;
use work.zpu_config.all;
use work.zpupkg.all;

entity Dhrystone_fast_ROM is
generic
	(
		maxAddrBitBRAM : integer := maxAddrBitBRAMLimit -- Specify your actual ROM size to save LEs and unnecessary block RAM usage.
	);
port (
	clk : in std_logic;
	areset : in std_logic := '0';
	from_zpu : in ZPU_ToROM;
	to_zpu : out ZPU_FromROM
);
end Dhrystone_fast_ROM;

architecture arch of Dhrystone_fast_ROM is

type ram_type is array(natural range 0 to ((2**(maxAddrBitBRAM+1))/4)-1) of std_logic_vector(wordSize-1 downto 0);

shared variable ram : ram_type :=
(
     0 => x"0b0b0b88",
     1 => x"dd040000",
     2 => x"00000000",
     3 => x"00000000",
     4 => x"00000000",
     5 => x"00000000",
     6 => x"00000000",
     7 => x"00000000",
     8 => x"88088c08",
     9 => x"90080b0b",
    10 => x"0b88e708",
    11 => x"2d900c8c",
    12 => x"0c880c04",
    13 => x"00000000",
    14 => x"00000000",
    15 => x"00000000",
    16 => x"71fd0608",
    17 => x"72830609",
    18 => x"81058205",
    19 => x"832b2a83",
    20 => x"ffff0652",
    21 => x"04000000",
    22 => x"00000000",
    23 => x"00000000",
    24 => x"71fd0608",
    25 => x"83ffff73",
    26 => x"83060981",
    27 => x"05820583",
    28 => x"2b2b0906",
    29 => x"7383ffff",
    30 => x"0b0b0b0b",
    31 => x"83a50400",
    32 => x"72098105",
    33 => x"72057373",
    34 => x"09060906",
    35 => x"73097306",
    36 => x"070a8106",
    37 => x"53510400",
    38 => x"00000000",
    39 => x"00000000",
    40 => x"72722473",
    41 => x"732e0753",
    42 => x"51040000",
    43 => x"00000000",
    44 => x"00000000",
    45 => x"00000000",
    46 => x"00000000",
    47 => x"00000000",
    48 => x"71737109",
    49 => x"71068106",
    50 => x"09810572",
    51 => x"0a100a72",
    52 => x"0a100a31",
    53 => x"050a8106",
    54 => x"51515351",
    55 => x"04000000",
    56 => x"72722673",
    57 => x"732e0753",
    58 => x"51040000",
    59 => x"00000000",
    60 => x"00000000",
    61 => x"00000000",
    62 => x"00000000",
    63 => x"00000000",
    64 => x"00000000",
    65 => x"00000000",
    66 => x"00000000",
    67 => x"00000000",
    68 => x"00000000",
    69 => x"00000000",
    70 => x"00000000",
    71 => x"00000000",
    72 => x"0b0b0b88",
    73 => x"ba040000",
    74 => x"00000000",
    75 => x"00000000",
    76 => x"00000000",
    77 => x"00000000",
    78 => x"00000000",
    79 => x"00000000",
    80 => x"720a722b",
    81 => x"0a535104",
    82 => x"00000000",
    83 => x"00000000",
    84 => x"00000000",
    85 => x"00000000",
    86 => x"00000000",
    87 => x"00000000",
    88 => x"72729f06",
    89 => x"0981050b",
    90 => x"0b0b889f",
    91 => x"05040000",
    92 => x"00000000",
    93 => x"00000000",
    94 => x"00000000",
    95 => x"00000000",
    96 => x"72722aff",
    97 => x"739f062a",
    98 => x"0974090a",
    99 => x"8106ff05",
   100 => x"06075351",
   101 => x"04000000",
   102 => x"00000000",
   103 => x"00000000",
   104 => x"71715351",
   105 => x"04067383",
   106 => x"06098105",
   107 => x"8205832b",
   108 => x"0b2b0772",
   109 => x"fc060c51",
   110 => x"51040000",
   111 => x"00000000",
   112 => x"72098105",
   113 => x"72050970",
   114 => x"81050906",
   115 => x"0a810653",
   116 => x"51040000",
   117 => x"00000000",
   118 => x"00000000",
   119 => x"00000000",
   120 => x"72098105",
   121 => x"72050970",
   122 => x"81050906",
   123 => x"0a098106",
   124 => x"53510400",
   125 => x"00000000",
   126 => x"00000000",
   127 => x"00000000",
   128 => x"71098105",
   129 => x"52040000",
   130 => x"00000000",
   131 => x"00000000",
   132 => x"00000000",
   133 => x"00000000",
   134 => x"00000000",
   135 => x"00000000",
   136 => x"72720981",
   137 => x"05055351",
   138 => x"04000000",
   139 => x"00000000",
   140 => x"00000000",
   141 => x"00000000",
   142 => x"00000000",
   143 => x"00000000",
   144 => x"72097206",
   145 => x"73730906",
   146 => x"07535104",
   147 => x"00000000",
   148 => x"00000000",
   149 => x"00000000",
   150 => x"00000000",
   151 => x"00000000",
   152 => x"71fc0608",
   153 => x"72830609",
   154 => x"81058305",
   155 => x"1010102a",
   156 => x"81ff0652",
   157 => x"04000000",
   158 => x"00000000",
   159 => x"00000000",
   160 => x"71fc0608",
   161 => x"0b0b0ba1",
   162 => x"ac738306",
   163 => x"10100508",
   164 => x"060b0b0b",
   165 => x"88a20400",
   166 => x"00000000",
   167 => x"00000000",
   168 => x"88088c08",
   169 => x"90087575",
   170 => x"0b0b0b9a",
   171 => x"9d2d5050",
   172 => x"88085690",
   173 => x"0c8c0c88",
   174 => x"0c510400",
   175 => x"00000000",
   176 => x"88088c08",
   177 => x"90087575",
   178 => x"0b0b0b9b",
   179 => x"cf2d5050",
   180 => x"88085690",
   181 => x"0c8c0c88",
   182 => x"0c510400",
   183 => x"00000000",
   184 => x"72097081",
   185 => x"0509060a",
   186 => x"8106ff05",
   187 => x"70547106",
   188 => x"73097274",
   189 => x"05ff0506",
   190 => x"07515151",
   191 => x"04000000",
   192 => x"72097081",
   193 => x"0509060a",
   194 => x"098106ff",
   195 => x"05705471",
   196 => x"06730972",
   197 => x"7405ff05",
   198 => x"06075151",
   199 => x"51040000",
   200 => x"05ff0504",
   201 => x"00000000",
   202 => x"00000000",
   203 => x"00000000",
   204 => x"00000000",
   205 => x"00000000",
   206 => x"00000000",
   207 => x"00000000",
   208 => x"04000000",
   209 => x"00000000",
   210 => x"00000000",
   211 => x"00000000",
   212 => x"00000000",
   213 => x"00000000",
   214 => x"00000000",
   215 => x"00000000",
   216 => x"71810552",
   217 => x"04000000",
   218 => x"00000000",
   219 => x"00000000",
   220 => x"00000000",
   221 => x"00000000",
   222 => x"00000000",
   223 => x"00000000",
   224 => x"00000000",
   225 => x"00000000",
   226 => x"00000000",
   227 => x"00000000",
   228 => x"00000000",
   229 => x"00000000",
   230 => x"00000000",
   231 => x"00000000",
   232 => x"02840572",
   233 => x"10100552",
   234 => x"04000000",
   235 => x"00000000",
   236 => x"00000000",
   237 => x"00000000",
   238 => x"00000000",
   239 => x"00000000",
   240 => x"00000000",
   241 => x"00000000",
   242 => x"00000000",
   243 => x"00000000",
   244 => x"00000000",
   245 => x"00000000",
   246 => x"00000000",
   247 => x"00000000",
   248 => x"717105ff",
   249 => x"05715351",
   250 => x"020d0400",
   251 => x"00000000",
   252 => x"00000000",
   253 => x"00000000",
   254 => x"00000000",
   255 => x"00000000",
   256 => x"10101010",
   257 => x"10101010",
   258 => x"10101010",
   259 => x"10101010",
   260 => x"10101010",
   261 => x"10101010",
   262 => x"10101010",
   263 => x"10101053",
   264 => x"51047381",
   265 => x"ff067383",
   266 => x"06098105",
   267 => x"83051010",
   268 => x"102b0772",
   269 => x"fc060c51",
   270 => x"51047272",
   271 => x"80728106",
   272 => x"ff050972",
   273 => x"06057110",
   274 => x"52720a10",
   275 => x"0a5372ed",
   276 => x"38515153",
   277 => x"51040000",
   278 => x"800488da",
   279 => x"0488da0b",
   280 => x"8fc10404",
   281 => x"00000000",
   282 => x"00046302",
   283 => x"c0050d02",
   284 => x"80c4050b",
   285 => x"0b0ba6d4",
   286 => x"5a5c807c",
   287 => x"7084055e",
   288 => x"08715f5f",
   289 => x"577d7084",
   290 => x"055f0856",
   291 => x"80587598",
   292 => x"2a76882b",
   293 => x"57557480",
   294 => x"2e82cd38",
   295 => x"7c802eb9",
   296 => x"38805d74",
   297 => x"80e42e81",
   298 => x"9f387480",
   299 => x"e42680dc",
   300 => x"387480e3",
   301 => x"2eba38a5",
   302 => x"518bf12d",
   303 => x"74518bf1",
   304 => x"2d821757",
   305 => x"81185883",
   306 => x"7825c338",
   307 => x"74ffb638",
   308 => x"7e880c02",
   309 => x"80c0050d",
   310 => x"0474a52e",
   311 => x"09810698",
   312 => x"38810b81",
   313 => x"19595d83",
   314 => x"7825ffa2",
   315 => x"3889cc04",
   316 => x"7b841d71",
   317 => x"08575d5a",
   318 => x"74518bf1",
   319 => x"2d811781",
   320 => x"19595783",
   321 => x"7825ff86",
   322 => x"3889cc04",
   323 => x"7480f32e",
   324 => x"098106ff",
   325 => x"a2387b84",
   326 => x"1d710870",
   327 => x"545b5d54",
   328 => x"8c922d80",
   329 => x"0bff1155",
   330 => x"53807325",
   331 => x"ff963878",
   332 => x"7081055a",
   333 => x"84e02d70",
   334 => x"52558bf1",
   335 => x"2d811774",
   336 => x"ff165654",
   337 => x"578aa904",
   338 => x"7b841d71",
   339 => x"080b0b0b",
   340 => x"a6d40b0b",
   341 => x"0b0ba684",
   342 => x"615f585e",
   343 => x"525d5372",
   344 => x"ba38b00b",
   345 => x"0b0b0ba6",
   346 => x"840b8580",
   347 => x"2d811454",
   348 => x"ff145473",
   349 => x"84e02d7b",
   350 => x"7081055d",
   351 => x"85802d81",
   352 => x"1a5a730b",
   353 => x"0b0ba684",
   354 => x"2e098106",
   355 => x"e338807b",
   356 => x"85802d79",
   357 => x"ff115553",
   358 => x"8aa9048a",
   359 => x"52725199",
   360 => x"f82d8808",
   361 => x"a1bc0584",
   362 => x"e02d7470",
   363 => x"81055685",
   364 => x"802d8a52",
   365 => x"725199d3",
   366 => x"2d880853",
   367 => x"8808dc38",
   368 => x"730b0b0b",
   369 => x"a6842ec6",
   370 => x"38ff1454",
   371 => x"7384e02d",
   372 => x"7b708105",
   373 => x"5d85802d",
   374 => x"811a5a73",
   375 => x"0b0b0ba6",
   376 => x"842effaa",
   377 => x"388af004",
   378 => x"76880c02",
   379 => x"80c0050d",
   380 => x"0402f805",
   381 => x"0d7352c0",
   382 => x"0870882a",
   383 => x"70810651",
   384 => x"51517080",
   385 => x"2ef13871",
   386 => x"c00c7188",
   387 => x"0c028805",
   388 => x"0d0402e8",
   389 => x"050d8078",
   390 => x"57557570",
   391 => x"84055708",
   392 => x"53805472",
   393 => x"982a7388",
   394 => x"2b545271",
   395 => x"802ea238",
   396 => x"c0087088",
   397 => x"2a708106",
   398 => x"51515170",
   399 => x"802ef138",
   400 => x"71c00c81",
   401 => x"15811555",
   402 => x"55837425",
   403 => x"d63871ca",
   404 => x"3874880c",
   405 => x"0298050d",
   406 => x"0402fc05",
   407 => x"0dc808f8",
   408 => x"80110888",
   409 => x"0c510284",
   410 => x"050d0402",
   411 => x"fc050d80",
   412 => x"c10b80f6",
   413 => x"a00b8580",
   414 => x"2d800b80",
   415 => x"f8b80c70",
   416 => x"880c0284",
   417 => x"050d0402",
   418 => x"f8050d80",
   419 => x"0b80f6a0",
   420 => x"0b84e02d",
   421 => x"52527080",
   422 => x"c12e9d38",
   423 => x"7180f8b8",
   424 => x"080780f8",
   425 => x"b80c80c2",
   426 => x"0b80f6a4",
   427 => x"0b85802d",
   428 => x"70880c02",
   429 => x"88050d04",
   430 => x"810b80f8",
   431 => x"b8080780",
   432 => x"f8b80c80",
   433 => x"c20b80f6",
   434 => x"a40b8580",
   435 => x"2d70880c",
   436 => x"0288050d",
   437 => x"0402f005",
   438 => x"0d757008",
   439 => x"8a055353",
   440 => x"80f6a00b",
   441 => x"84e02d51",
   442 => x"7080c12e",
   443 => x"8c3873f0",
   444 => x"3870880c",
   445 => x"0290050d",
   446 => x"04ff1270",
   447 => x"80f69c08",
   448 => x"31740c88",
   449 => x"0c029005",
   450 => x"0d0402ec",
   451 => x"050d80f6",
   452 => x"c8085574",
   453 => x"802e8c38",
   454 => x"76750871",
   455 => x"0c80f6c8",
   456 => x"0856548c",
   457 => x"155380f6",
   458 => x"9c08528a",
   459 => x"5197a92d",
   460 => x"73880c02",
   461 => x"94050d04",
   462 => x"02e8050d",
   463 => x"77700856",
   464 => x"56b05380",
   465 => x"f6c80852",
   466 => x"74519efb",
   467 => x"2d850b8c",
   468 => x"170c850b",
   469 => x"8c160c75",
   470 => x"08750c80",
   471 => x"f6c80854",
   472 => x"73802e8a",
   473 => x"38730875",
   474 => x"0c80f6c8",
   475 => x"08548c14",
   476 => x"5380f69c",
   477 => x"08528a51",
   478 => x"97a92d84",
   479 => x"1508ae38",
   480 => x"860b8c16",
   481 => x"0c881552",
   482 => x"88160851",
   483 => x"96c32d80",
   484 => x"f6c80870",
   485 => x"08760c54",
   486 => x"8c157054",
   487 => x"548a5273",
   488 => x"085197a9",
   489 => x"2d73880c",
   490 => x"0298050d",
   491 => x"04750854",
   492 => x"b0537352",
   493 => x"75519efb",
   494 => x"2d73880c",
   495 => x"0298050d",
   496 => x"0402c805",
   497 => x"0d80f5b4",
   498 => x"0b80f5e8",
   499 => x"0c80f5ec",
   500 => x"0b80f6c8",
   501 => x"0c80f5b4",
   502 => x"0b80f5ec",
   503 => x"0c800b80",
   504 => x"f5ec0b84",
   505 => x"050c820b",
   506 => x"80f5ec0b",
   507 => x"88050ca8",
   508 => x"0b80f5ec",
   509 => x"0b8c050c",
   510 => x"9f53a1d0",
   511 => x"5280f5fc",
   512 => x"519efb2d",
   513 => x"9f53a1f0",
   514 => x"5280f898",
   515 => x"519efb2d",
   516 => x"8a0bb480",
   517 => x"0ca4d051",
   518 => x"88eb2da2",
   519 => x"905188eb",
   520 => x"2da4d051",
   521 => x"88eb2da6",
   522 => x"8008802e",
   523 => x"849b38a2",
   524 => x"c05188eb",
   525 => x"2da4d051",
   526 => x"88eb2da5",
   527 => x"fc0852a2",
   528 => x"ec5188eb",
   529 => x"2dc808f8",
   530 => x"80110870",
   531 => x"a7a00c57",
   532 => x"55815880",
   533 => x"0ba5fc08",
   534 => x"2582dc38",
   535 => x"02ac055b",
   536 => x"80c10b80",
   537 => x"f6a00b85",
   538 => x"802d810b",
   539 => x"80f8b80c",
   540 => x"80c20b80",
   541 => x"f6a40b85",
   542 => x"802d825c",
   543 => x"835a9f53",
   544 => x"a39c5280",
   545 => x"f6a8519e",
   546 => x"fb2d815d",
   547 => x"800b80f6",
   548 => x"a85380f8",
   549 => x"98525598",
   550 => x"db2d8808",
   551 => x"752e0981",
   552 => x"06833881",
   553 => x"557480f8",
   554 => x"b80c7b70",
   555 => x"57557483",
   556 => x"25a13874",
   557 => x"101015fd",
   558 => x"055e02b8",
   559 => x"05fc0553",
   560 => x"83527551",
   561 => x"97a92d81",
   562 => x"1c705d70",
   563 => x"57558375",
   564 => x"24e1387d",
   565 => x"547453a7",
   566 => x"a45280f6",
   567 => x"d05197bb",
   568 => x"2d80f6c8",
   569 => x"08700857",
   570 => x"57b05376",
   571 => x"5275519e",
   572 => x"fb2d850b",
   573 => x"8c180c85",
   574 => x"0b8c170c",
   575 => x"7608760c",
   576 => x"80f6c808",
   577 => x"5574802e",
   578 => x"8a387408",
   579 => x"760c80f6",
   580 => x"c808558c",
   581 => x"155380f6",
   582 => x"9c08528a",
   583 => x"5197a92d",
   584 => x"84160883",
   585 => x"dd38860b",
   586 => x"8c170c88",
   587 => x"16528817",
   588 => x"085196c3",
   589 => x"2d80f6c8",
   590 => x"08700877",
   591 => x"0c558c16",
   592 => x"7054578a",
   593 => x"52760851",
   594 => x"97a92d80",
   595 => x"c10b80f6",
   596 => x"a40b84e0",
   597 => x"2d565675",
   598 => x"7526a538",
   599 => x"80c35275",
   600 => x"5198a72d",
   601 => x"88087d2e",
   602 => x"82e73881",
   603 => x"167081ff",
   604 => x"0680f6a4",
   605 => x"0b84e02d",
   606 => x"57575774",
   607 => x"7627dd38",
   608 => x"797c297e",
   609 => x"53519a9d",
   610 => x"2d88085c",
   611 => x"88088a05",
   612 => x"80f6a00b",
   613 => x"84e02d80",
   614 => x"f69c0859",
   615 => x"57557580",
   616 => x"c12e82f9",
   617 => x"3878f738",
   618 => x"811858a5",
   619 => x"fc087825",
   620 => x"fdae38a7",
   621 => x"a00856c8",
   622 => x"08f88011",
   623 => x"087080f5",
   624 => x"e40c7078",
   625 => x"3170a79c",
   626 => x"0c54a3bc",
   627 => x"535c5a88",
   628 => x"eb2da79c",
   629 => x"085680f7",
   630 => x"762580f3",
   631 => x"38a5fc08",
   632 => x"70537687",
   633 => x"e8295257",
   634 => x"9a9d2d88",
   635 => x"08a7940c",
   636 => x"75527687",
   637 => x"e829519a",
   638 => x"9d2d8808",
   639 => x"a7980c75",
   640 => x"527684b9",
   641 => x"29519a9d",
   642 => x"2d880880",
   643 => x"f6cc0ca3",
   644 => x"cc5188eb",
   645 => x"2da79408",
   646 => x"52a3fc51",
   647 => x"88eb2da4",
   648 => x"845188eb",
   649 => x"2da79808",
   650 => x"52a3fc51",
   651 => x"88eb2d80",
   652 => x"f6cc0852",
   653 => x"a4b45188",
   654 => x"eb2da4d0",
   655 => x"5188eb2d",
   656 => x"800b880c",
   657 => x"02b8050d",
   658 => x"04a4d451",
   659 => x"90b204a5",
   660 => x"845188eb",
   661 => x"2da5bc51",
   662 => x"88eb2da4",
   663 => x"d05188eb",
   664 => x"2da79c08",
   665 => x"a5fc0870",
   666 => x"547187e8",
   667 => x"29535856",
   668 => x"9a9d2d88",
   669 => x"08a7940c",
   670 => x"75527687",
   671 => x"e829519a",
   672 => x"9d2d8808",
   673 => x"a7980c75",
   674 => x"527684b9",
   675 => x"29519a9d",
   676 => x"2d880880",
   677 => x"f6cc0ca3",
   678 => x"cc5188eb",
   679 => x"2da79408",
   680 => x"52a3fc51",
   681 => x"88eb2da4",
   682 => x"845188eb",
   683 => x"2da79808",
   684 => x"52a3fc51",
   685 => x"88eb2d80",
   686 => x"f6cc0852",
   687 => x"a4b45188",
   688 => x"eb2da4d0",
   689 => x"5188eb2d",
   690 => x"800b880c",
   691 => x"02b8050d",
   692 => x"0402b805",
   693 => x"f8055280",
   694 => x"5196c32d",
   695 => x"9f53a5dc",
   696 => x"5280f6a8",
   697 => x"519efb2d",
   698 => x"777880f6",
   699 => x"9c0c8117",
   700 => x"7081ff06",
   701 => x"80f6a40b",
   702 => x"84e02d58",
   703 => x"58585a92",
   704 => x"fb047608",
   705 => x"56b05375",
   706 => x"5276519e",
   707 => x"fb2d80c1",
   708 => x"0b80f6a4",
   709 => x"0b84e02d",
   710 => x"565692d7",
   711 => x"04ff1570",
   712 => x"78317c0c",
   713 => x"59805993",
   714 => x"a80402f8",
   715 => x"050d7382",
   716 => x"32700981",
   717 => x"05707207",
   718 => x"8025880c",
   719 => x"52520288",
   720 => x"050d0402",
   721 => x"f4050d74",
   722 => x"76715354",
   723 => x"5271822e",
   724 => x"83388351",
   725 => x"71812e9b",
   726 => x"38817226",
   727 => x"a0387182",
   728 => x"2ebc3871",
   729 => x"842eac38",
   730 => x"70730c70",
   731 => x"880c028c",
   732 => x"050d0480",
   733 => x"e40b80f6",
   734 => x"9c08258c",
   735 => x"3880730c",
   736 => x"70880c02",
   737 => x"8c050d04",
   738 => x"83730c70",
   739 => x"880c028c",
   740 => x"050d0482",
   741 => x"730c7088",
   742 => x"0c028c05",
   743 => x"0d048173",
   744 => x"0c70880c",
   745 => x"028c050d",
   746 => x"0402fc05",
   747 => x"0d747414",
   748 => x"8205710c",
   749 => x"880c0284",
   750 => x"050d0402",
   751 => x"d8050d7b",
   752 => x"7d7f6185",
   753 => x"1270822b",
   754 => x"75117074",
   755 => x"71708405",
   756 => x"530c5a5a",
   757 => x"5d5b760c",
   758 => x"7980f818",
   759 => x"0c798612",
   760 => x"5257585a",
   761 => x"5a767624",
   762 => x"993876b3",
   763 => x"29822b79",
   764 => x"11515376",
   765 => x"73708405",
   766 => x"550c8114",
   767 => x"54757425",
   768 => x"f2387681",
   769 => x"cc2919fc",
   770 => x"11088105",
   771 => x"fc120c7a",
   772 => x"1970089f",
   773 => x"a0130c58",
   774 => x"56850b80",
   775 => x"f69c0c75",
   776 => x"880c02a8",
   777 => x"050d0402",
   778 => x"f4050d02",
   779 => x"930584e0",
   780 => x"2d518002",
   781 => x"84059705",
   782 => x"84e02d54",
   783 => x"5270732e",
   784 => x"89387188",
   785 => x"0c028c05",
   786 => x"0d047080",
   787 => x"f6a00b85",
   788 => x"802d810b",
   789 => x"880c028c",
   790 => x"050d0402",
   791 => x"dc050d7a",
   792 => x"7c595682",
   793 => x"0b831955",
   794 => x"55741670",
   795 => x"84e02d75",
   796 => x"84e02d5b",
   797 => x"51537279",
   798 => x"2e80c738",
   799 => x"80c10b81",
   800 => x"16811656",
   801 => x"56578275",
   802 => x"25df38ff",
   803 => x"a9177081",
   804 => x"ff065559",
   805 => x"73822683",
   806 => x"38875581",
   807 => x"537680d2",
   808 => x"2e983877",
   809 => x"527551a0",
   810 => x"942d8053",
   811 => x"72880825",
   812 => x"89388715",
   813 => x"80f69c0c",
   814 => x"81537288",
   815 => x"0c02a405",
   816 => x"0d047280",
   817 => x"f6a00b85",
   818 => x"802d8275",
   819 => x"25ff9a38",
   820 => x"998b0494",
   821 => x"0802940c",
   822 => x"fd3d0d80",
   823 => x"5394088c",
   824 => x"05085294",
   825 => x"08880508",
   826 => x"5182de3f",
   827 => x"88087088",
   828 => x"0c54853d",
   829 => x"0d940c04",
   830 => x"94080294",
   831 => x"0cfd3d0d",
   832 => x"81539408",
   833 => x"8c050852",
   834 => x"94088805",
   835 => x"085182b9",
   836 => x"3f880870",
   837 => x"880c5485",
   838 => x"3d0d940c",
   839 => x"04940802",
   840 => x"940cf93d",
   841 => x"0d800b94",
   842 => x"08fc050c",
   843 => x"94088805",
   844 => x"088025ab",
   845 => x"38940888",
   846 => x"05083094",
   847 => x"0888050c",
   848 => x"800b9408",
   849 => x"f4050c94",
   850 => x"08fc0508",
   851 => x"8838810b",
   852 => x"9408f405",
   853 => x"0c9408f4",
   854 => x"05089408",
   855 => x"fc050c94",
   856 => x"088c0508",
   857 => x"8025ab38",
   858 => x"94088c05",
   859 => x"08309408",
   860 => x"8c050c80",
   861 => x"0b9408f0",
   862 => x"050c9408",
   863 => x"fc050888",
   864 => x"38810b94",
   865 => x"08f0050c",
   866 => x"9408f005",
   867 => x"089408fc",
   868 => x"050c8053",
   869 => x"94088c05",
   870 => x"08529408",
   871 => x"88050851",
   872 => x"81a73f88",
   873 => x"08709408",
   874 => x"f8050c54",
   875 => x"9408fc05",
   876 => x"08802e8c",
   877 => x"389408f8",
   878 => x"05083094",
   879 => x"08f8050c",
   880 => x"9408f805",
   881 => x"0870880c",
   882 => x"54893d0d",
   883 => x"940c0494",
   884 => x"0802940c",
   885 => x"fb3d0d80",
   886 => x"0b9408fc",
   887 => x"050c9408",
   888 => x"88050880",
   889 => x"25933894",
   890 => x"08880508",
   891 => x"30940888",
   892 => x"050c810b",
   893 => x"9408fc05",
   894 => x"0c94088c",
   895 => x"05088025",
   896 => x"8c389408",
   897 => x"8c050830",
   898 => x"94088c05",
   899 => x"0c815394",
   900 => x"088c0508",
   901 => x"52940888",
   902 => x"050851ad",
   903 => x"3f880870",
   904 => x"9408f805",
   905 => x"0c549408",
   906 => x"fc050880",
   907 => x"2e8c3894",
   908 => x"08f80508",
   909 => x"309408f8",
   910 => x"050c9408",
   911 => x"f8050870",
   912 => x"880c5487",
   913 => x"3d0d940c",
   914 => x"04940802",
   915 => x"940cfd3d",
   916 => x"0d810b94",
   917 => x"08fc050c",
   918 => x"800b9408",
   919 => x"f8050c94",
   920 => x"088c0508",
   921 => x"94088805",
   922 => x"0827ac38",
   923 => x"9408fc05",
   924 => x"08802ea3",
   925 => x"38800b94",
   926 => x"088c0508",
   927 => x"24993894",
   928 => x"088c0508",
   929 => x"1094088c",
   930 => x"050c9408",
   931 => x"fc050810",
   932 => x"9408fc05",
   933 => x"0cc93994",
   934 => x"08fc0508",
   935 => x"802e80c9",
   936 => x"3894088c",
   937 => x"05089408",
   938 => x"88050826",
   939 => x"a1389408",
   940 => x"88050894",
   941 => x"088c0508",
   942 => x"31940888",
   943 => x"050c9408",
   944 => x"f8050894",
   945 => x"08fc0508",
   946 => x"079408f8",
   947 => x"050c9408",
   948 => x"fc050881",
   949 => x"2a9408fc",
   950 => x"050c9408",
   951 => x"8c050881",
   952 => x"2a94088c",
   953 => x"050cffaf",
   954 => x"39940890",
   955 => x"0508802e",
   956 => x"8f389408",
   957 => x"88050870",
   958 => x"9408f405",
   959 => x"0c518d39",
   960 => x"9408f805",
   961 => x"08709408",
   962 => x"f4050c51",
   963 => x"9408f405",
   964 => x"08880c85",
   965 => x"3d0d940c",
   966 => x"04940802",
   967 => x"940cff3d",
   968 => x"0d800b94",
   969 => x"08fc050c",
   970 => x"94088805",
   971 => x"088106ff",
   972 => x"11700970",
   973 => x"94088c05",
   974 => x"08069408",
   975 => x"fc050811",
   976 => x"9408fc05",
   977 => x"0c940888",
   978 => x"0508812a",
   979 => x"94088805",
   980 => x"0c94088c",
   981 => x"05081094",
   982 => x"088c050c",
   983 => x"51515151",
   984 => x"94088805",
   985 => x"08802e84",
   986 => x"38ffbd39",
   987 => x"9408fc05",
   988 => x"0870880c",
   989 => x"51833d0d",
   990 => x"940c04fc",
   991 => x"3d0d7670",
   992 => x"797b5555",
   993 => x"55558f72",
   994 => x"278c3872",
   995 => x"75078306",
   996 => x"5170802e",
   997 => x"a738ff12",
   998 => x"5271ff2e",
   999 => x"98387270",
  1000 => x"81055433",
  1001 => x"74708105",
  1002 => x"5634ff12",
  1003 => x"5271ff2e",
  1004 => x"098106ea",
  1005 => x"3874880c",
  1006 => x"863d0d04",
  1007 => x"74517270",
  1008 => x"84055408",
  1009 => x"71708405",
  1010 => x"530c7270",
  1011 => x"84055408",
  1012 => x"71708405",
  1013 => x"530c7270",
  1014 => x"84055408",
  1015 => x"71708405",
  1016 => x"530c7270",
  1017 => x"84055408",
  1018 => x"71708405",
  1019 => x"530cf012",
  1020 => x"52718f26",
  1021 => x"c9388372",
  1022 => x"27953872",
  1023 => x"70840554",
  1024 => x"08717084",
  1025 => x"05530cfc",
  1026 => x"12527183",
  1027 => x"26ed3870",
  1028 => x"54ff8339",
  1029 => x"fb3d0d77",
  1030 => x"79707207",
  1031 => x"83065354",
  1032 => x"52709338",
  1033 => x"71737308",
  1034 => x"54565471",
  1035 => x"73082e80",
  1036 => x"c4387375",
  1037 => x"54527133",
  1038 => x"7081ff06",
  1039 => x"52547080",
  1040 => x"2e9d3872",
  1041 => x"33557075",
  1042 => x"2e098106",
  1043 => x"95388112",
  1044 => x"81147133",
  1045 => x"7081ff06",
  1046 => x"54565452",
  1047 => x"70e53872",
  1048 => x"33557381",
  1049 => x"ff067581",
  1050 => x"ff067171",
  1051 => x"31880c52",
  1052 => x"52873d0d",
  1053 => x"04710970",
  1054 => x"f7fbfdff",
  1055 => x"140670f8",
  1056 => x"84828180",
  1057 => x"06515151",
  1058 => x"70973884",
  1059 => x"14841671",
  1060 => x"08545654",
  1061 => x"7175082e",
  1062 => x"dc387375",
  1063 => x"5452ff96",
  1064 => x"39800b88",
  1065 => x"0c873d0d",
  1066 => x"04000000",
  1067 => x"00ffffff",
  1068 => x"ff00ffff",
  1069 => x"ffff00ff",
  1070 => x"ffffff00",
  1071 => x"30313233",
  1072 => x"34353637",
  1073 => x"38394142",
  1074 => x"43444546",
  1075 => x"00000000",
  1076 => x"44485259",
  1077 => x"53544f4e",
  1078 => x"45205052",
  1079 => x"4f475241",
  1080 => x"4d2c2053",
  1081 => x"4f4d4520",
  1082 => x"53545249",
  1083 => x"4e470000",
  1084 => x"44485259",
  1085 => x"53544f4e",
  1086 => x"45205052",
  1087 => x"4f475241",
  1088 => x"4d2c2031",
  1089 => x"27535420",
  1090 => x"53545249",
  1091 => x"4e470000",
  1092 => x"44687279",
  1093 => x"73746f6e",
  1094 => x"65204265",
  1095 => x"6e63686d",
  1096 => x"61726b2c",
  1097 => x"20566572",
  1098 => x"73696f6e",
  1099 => x"20322e31",
  1100 => x"20284c61",
  1101 => x"6e677561",
  1102 => x"67653a20",
  1103 => x"43290a00",
  1104 => x"50726f67",
  1105 => x"72616d20",
  1106 => x"636f6d70",
  1107 => x"696c6564",
  1108 => x"20776974",
  1109 => x"68202772",
  1110 => x"65676973",
  1111 => x"74657227",
  1112 => x"20617474",
  1113 => x"72696275",
  1114 => x"74650a00",
  1115 => x"45786563",
  1116 => x"7574696f",
  1117 => x"6e207374",
  1118 => x"61727473",
  1119 => x"2c202564",
  1120 => x"2072756e",
  1121 => x"73207468",
  1122 => x"726f7567",
  1123 => x"68204468",
  1124 => x"72797374",
  1125 => x"6f6e650a",
  1126 => x"00000000",
  1127 => x"44485259",
  1128 => x"53544f4e",
  1129 => x"45205052",
  1130 => x"4f475241",
  1131 => x"4d2c2032",
  1132 => x"274e4420",
  1133 => x"53545249",
  1134 => x"4e470000",
  1135 => x"55736572",
  1136 => x"2074696d",
  1137 => x"653a2025",
  1138 => x"640a0000",
  1139 => x"4d696372",
  1140 => x"6f736563",
  1141 => x"6f6e6473",
  1142 => x"20666f72",
  1143 => x"206f6e65",
  1144 => x"2072756e",
  1145 => x"20746872",
  1146 => x"6f756768",
  1147 => x"20446872",
  1148 => x"7973746f",
  1149 => x"6e653a20",
  1150 => x"00000000",
  1151 => x"2564200a",
  1152 => x"00000000",
  1153 => x"44687279",
  1154 => x"73746f6e",
  1155 => x"65732070",
  1156 => x"65722053",
  1157 => x"65636f6e",
  1158 => x"643a2020",
  1159 => x"20202020",
  1160 => x"20202020",
  1161 => x"20202020",
  1162 => x"20202020",
  1163 => x"20202020",
  1164 => x"00000000",
  1165 => x"56415820",
  1166 => x"4d495053",
  1167 => x"20726174",
  1168 => x"696e6720",
  1169 => x"2a203130",
  1170 => x"3030203d",
  1171 => x"20256420",
  1172 => x"0a000000",
  1173 => x"50726f67",
  1174 => x"72616d20",
  1175 => x"636f6d70",
  1176 => x"696c6564",
  1177 => x"20776974",
  1178 => x"686f7574",
  1179 => x"20277265",
  1180 => x"67697374",
  1181 => x"65722720",
  1182 => x"61747472",
  1183 => x"69627574",
  1184 => x"650a0000",
  1185 => x"4d656173",
  1186 => x"75726564",
  1187 => x"2074696d",
  1188 => x"6520746f",
  1189 => x"6f20736d",
  1190 => x"616c6c20",
  1191 => x"746f206f",
  1192 => x"62746169",
  1193 => x"6e206d65",
  1194 => x"616e696e",
  1195 => x"6766756c",
  1196 => x"20726573",
  1197 => x"756c7473",
  1198 => x"0a000000",
  1199 => x"506c6561",
  1200 => x"73652069",
  1201 => x"6e637265",
  1202 => x"61736520",
  1203 => x"6e756d62",
  1204 => x"6572206f",
  1205 => x"66207275",
  1206 => x"6e730a00",
  1207 => x"44485259",
  1208 => x"53544f4e",
  1209 => x"45205052",
  1210 => x"4f475241",
  1211 => x"4d2c2033",
  1212 => x"27524420",
  1213 => x"53545249",
  1214 => x"4e470000",
  1215 => x"000061a8",
  1216 => x"00000000",
	others => x"00000000"
);

begin

process (clk)
begin
	if (clk'event and clk = '1') then
		if (from_zpu.memAWriteEnable = '1') and (from_zpu.memBWriteEnable = '1') and (from_zpu.memAAddr=from_zpu.memBAddr) and (from_zpu.memAWrite/=from_zpu.memBWrite) then
			report "write collision" severity failure;
		end if;
	
		if (from_zpu.memAWriteEnable = '1') then
			ram(to_integer(unsigned(from_zpu.memAAddr(maxAddrBitBRAM downto 2)))) := from_zpu.memAWrite;
			to_zpu.memARead <= from_zpu.memAWrite;
		else
			to_zpu.memARead <= ram(to_integer(unsigned(from_zpu.memAAddr(maxAddrBitBRAM downto 2))));
		end if;
	end if;
end process;

process (clk)
begin
	if (clk'event and clk = '1') then
		if (from_zpu.memBWriteEnable = '1') then
			ram(to_integer(unsigned(from_zpu.memBAddr(maxAddrBitBRAM downto 2)))) := from_zpu.memBWrite;
			to_zpu.memBRead <= from_zpu.memBWrite;
		else
			to_zpu.memBRead <= ram(to_integer(unsigned(from_zpu.memBAddr(maxAddrBitBRAM downto 2))));
		end if;
	end if;
end process;


end arch;

