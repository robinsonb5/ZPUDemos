-- ZPU
--
-- Copyright 2004-2008 oharboe - �yvind Harboe - oyvind.harboe@zylin.com
-- Modified by Alastair M. Robinson for the ZPUFlex project.
--
-- The FreeBSD license
-- 
-- Redistribution and use in source and binary forms, with or without
-- modification, are permitted provided that the following conditions
-- are met:
-- 
-- 1. Redistributions of source code must retain the above copyright
--    notice, this list of conditions and the following disclaimer.
-- 2. Redistributions in binary form must reproduce the above
--    copyright notice, this list of conditions and the following
--    disclaimer in the documentation and/or other materials
--    provided with the distribution.
-- 
-- THIS SOFTWARE IS PROVIDED BY THE ZPU PROJECT ``AS IS'' AND ANY
-- EXPRESS OR IMPLIED WARRANTIES, INCLUDING, BUT NOT LIMITED TO,
-- THE IMPLIED WARRANTIES OF MERCHANTABILITY AND FITNESS FOR A
-- PARTICULAR PURPOSE ARE DISCLAIMED. IN NO EVENT SHALL THE
-- ZPU PROJECT OR CONTRIBUTORS BE LIABLE FOR ANY DIRECT,
-- INDIRECT, INCIDENTAL, SPECIAL, EXEMPLARY, OR CONSEQUENTIAL DAMAGES
-- (INCLUDING, BUT NOT LIMITED TO, PROCUREMENT OF SUBSTITUTE GOODS
-- OR SERVICES; LOSS OF USE, DATA, OR PROFITS; OR BUSINESS INTERRUPTION)
-- HOWEVER CAUSED AND ON ANY THEORY OF LIABILITY, WHETHER IN CONTRACT,
-- STRICT LIABILITY, OR TORT (INCLUDING NEGLIGENCE OR OTHERWISE)
-- ARISING IN ANY WAY OUT OF THE USE OF THIS SOFTWARE, EVEN IF
-- ADVISED OF THE POSSIBILITY OF SUCH DAMAGE.
-- 
-- The views and conclusions contained in the software and documentation
-- are those of the authors and should not be interpreted as representing
-- official policies, either expressed or implied, of the ZPU Project.

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;


library work;
use work.zpupkg.all;

entity SDRAMTest_ROM is
generic
	(
		maxAddrBitBRAM : integer := maxAddrBitBRAMLimit -- Specify your actual ROM size to save LEs and unnecessary block RAM usage.
	);
port (
	clk : in std_logic;
	areset : in std_logic := '0';
	from_zpu : in ZPU_ToROM;
	to_zpu : out ZPU_FromROM
);
end SDRAMTest_ROM;

architecture arch of SDRAMTest_ROM is

type ram_type is array(natural range 0 to ((2**(maxAddrBitBRAM+1))/4)-1) of std_logic_vector(wordSize-1 downto 0);

shared variable ram : ram_type :=
(
     0 => x"84808080",
     1 => x"8c0b8480",
     2 => x"8081e004",
     3 => x"00848080",
     4 => x"808c04ff",
     5 => x"0d800404",
     6 => x"40000017",
     7 => x"00000000",
     8 => x"848080a8",
     9 => x"c4088480",
    10 => x"80a8c808",
    11 => x"848080a8",
    12 => x"cc088480",
    13 => x"80809808",
    14 => x"2d848080",
    15 => x"a8cc0c84",
    16 => x"8080a8c8",
    17 => x"0c848080",
    18 => x"a8c40c04",
    19 => x"00000000",
    20 => x"00000000",
    21 => x"00000000",
    22 => x"00000000",
    23 => x"00000000",
    24 => x"71fd0608",
    25 => x"72830609",
    26 => x"81058205",
    27 => x"832b2a83",
    28 => x"ffff0652",
    29 => x"0471fc06",
    30 => x"08728306",
    31 => x"09810583",
    32 => x"05101010",
    33 => x"2a81ff06",
    34 => x"520471fd",
    35 => x"060883ff",
    36 => x"ff738306",
    37 => x"09810582",
    38 => x"05832b2b",
    39 => x"09067383",
    40 => x"ffff0673",
    41 => x"83060981",
    42 => x"05820583",
    43 => x"2b0b2b07",
    44 => x"72fc060c",
    45 => x"51510471",
    46 => x"fc060884",
    47 => x"808099e0",
    48 => x"73830610",
    49 => x"10050806",
    50 => x"7381ff06",
    51 => x"73830609",
    52 => x"81058305",
    53 => x"1010102b",
    54 => x"0772fc06",
    55 => x"0c515104",
    56 => x"848080a8",
    57 => x"c4708480",
    58 => x"80a9e427",
    59 => x"8e388071",
    60 => x"70840553",
    61 => x"0c848080",
    62 => x"81e50484",
    63 => x"8080808c",
    64 => x"51848080",
    65 => x"95fc0402",
    66 => x"c0050d02",
    67 => x"80c4055b",
    68 => x"80707c70",
    69 => x"84055e08",
    70 => x"725f5f5f",
    71 => x"5a7c7084",
    72 => x"055e0857",
    73 => x"80597698",
    74 => x"2a77882b",
    75 => x"58557480",
    76 => x"2e82e738",
    77 => x"7b802e80",
    78 => x"d338805c",
    79 => x"7480e42e",
    80 => x"81d83874",
    81 => x"80f82e81",
    82 => x"d1387480",
    83 => x"e42e81dc",
    84 => x"387480e4",
    85 => x"2680f138",
    86 => x"7480e32e",
    87 => x"80c838a5",
    88 => x"51848080",
    89 => x"85db2d74",
    90 => x"51848080",
    91 => x"85db2d82",
    92 => x"1a811a5a",
    93 => x"5a837925",
    94 => x"ffac3874",
    95 => x"ff9f387e",
    96 => x"848080a8",
    97 => x"c40c0280",
    98 => x"c0050d04",
    99 => x"74a52e09",
   100 => x"81069b38",
   101 => x"810b811a",
   102 => x"5a5c8379",
   103 => x"25ff8738",
   104 => x"84808082",
   105 => x"fb047a84",
   106 => x"1c710857",
   107 => x"5c547451",
   108 => x"84808085",
   109 => x"db2d811a",
   110 => x"811a5a5a",
   111 => x"837925fe",
   112 => x"e5388480",
   113 => x"8082fb04",
   114 => x"7480f32e",
   115 => x"81d93874",
   116 => x"80f82e09",
   117 => x"8106ff87",
   118 => x"387d5380",
   119 => x"587d782e",
   120 => x"81e23887",
   121 => x"56729c2a",
   122 => x"73842b54",
   123 => x"5271802e",
   124 => x"83388158",
   125 => x"b7125471",
   126 => x"89248438",
   127 => x"b0125477",
   128 => x"80ea38ff",
   129 => x"16567580",
   130 => x"25db3881",
   131 => x"19598379",
   132 => x"25fe9338",
   133 => x"84808082",
   134 => x"fb047a84",
   135 => x"1c710840",
   136 => x"5c527480",
   137 => x"e42e0981",
   138 => x"06fea638",
   139 => x"7d538058",
   140 => x"7d782e81",
   141 => x"8f388756",
   142 => x"729c2a73",
   143 => x"842b5452",
   144 => x"71802e83",
   145 => x"388158b7",
   146 => x"12547189",
   147 => x"248438b0",
   148 => x"125477af",
   149 => x"38ff1656",
   150 => x"758025dc",
   151 => x"38811959",
   152 => x"837925fd",
   153 => x"c1388480",
   154 => x"8082fb04",
   155 => x"73518480",
   156 => x"8085db2d",
   157 => x"ff165675",
   158 => x"8025fee9",
   159 => x"38848080",
   160 => x"848b0473",
   161 => x"51848080",
   162 => x"85db2dff",
   163 => x"16567580",
   164 => x"25ffa538",
   165 => x"84808084",
   166 => x"dd047984",
   167 => x"8080a8c4",
   168 => x"0c0280c0",
   169 => x"050d047a",
   170 => x"841c7108",
   171 => x"535c5384",
   172 => x"80808680",
   173 => x"2d811959",
   174 => x"837925fc",
   175 => x"e9388480",
   176 => x"8082fb04",
   177 => x"b0518480",
   178 => x"8085db2d",
   179 => x"81195983",
   180 => x"7925fcd2",
   181 => x"38848080",
   182 => x"82fb0402",
   183 => x"f8050d73",
   184 => x"52c00870",
   185 => x"882a7081",
   186 => x"06515151",
   187 => x"70802ef1",
   188 => x"3871c00c",
   189 => x"71848080",
   190 => x"a8c40c02",
   191 => x"88050d04",
   192 => x"02e8050d",
   193 => x"80785755",
   194 => x"75708405",
   195 => x"57085380",
   196 => x"5472982a",
   197 => x"73882b54",
   198 => x"5271802e",
   199 => x"a238c008",
   200 => x"70882a70",
   201 => x"81065151",
   202 => x"5170802e",
   203 => x"f13871c0",
   204 => x"0c811581",
   205 => x"15555583",
   206 => x"7425d638",
   207 => x"71ca3874",
   208 => x"848080a8",
   209 => x"c40c0298",
   210 => x"050d0402",
   211 => x"f4050d74",
   212 => x"76525380",
   213 => x"71259038",
   214 => x"70527270",
   215 => x"84055408",
   216 => x"ff135351",
   217 => x"71f43802",
   218 => x"8c050d04",
   219 => x"02d4050d",
   220 => x"7c7e5c58",
   221 => x"810b8480",
   222 => x"8099f058",
   223 => x"5a835976",
   224 => x"08780c77",
   225 => x"08770856",
   226 => x"5473752e",
   227 => x"94387708",
   228 => x"53745284",
   229 => x"80809a80",
   230 => x"51848080",
   231 => x"82872d80",
   232 => x"5a775680",
   233 => x"7b259038",
   234 => x"7a557570",
   235 => x"84055708",
   236 => x"ff165654",
   237 => x"74f43877",
   238 => x"08770856",
   239 => x"5675752e",
   240 => x"94387708",
   241 => x"53745284",
   242 => x"80809ac0",
   243 => x"51848080",
   244 => x"82872d80",
   245 => x"5aff1984",
   246 => x"18585978",
   247 => x"8025ff9f",
   248 => x"38798480",
   249 => x"80a8c40c",
   250 => x"02ac050d",
   251 => x"0402e405",
   252 => x"0d787a55",
   253 => x"56817608",
   254 => x"84180888",
   255 => x"19088c1a",
   256 => x"08515151",
   257 => x"545785aa",
   258 => x"d5aad576",
   259 => x"0cfad5aa",
   260 => x"d5aa0b8c",
   261 => x"170ccc76",
   262 => x"34b30b8f",
   263 => x"17347508",
   264 => x"5372fce2",
   265 => x"d5aad52e",
   266 => x"92387508",
   267 => x"52848080",
   268 => x"9b805184",
   269 => x"80808287",
   270 => x"2d80578c",
   271 => x"16085574",
   272 => x"fad5aad4",
   273 => x"b32e9338",
   274 => x"8c160852",
   275 => x"8480809b",
   276 => x"bc518480",
   277 => x"8082872d",
   278 => x"8057920b",
   279 => x"811734fd",
   280 => x"dc0b8e17",
   281 => x"23750853",
   282 => x"72fce0c9",
   283 => x"aad52e92",
   284 => x"38750852",
   285 => x"8480809b",
   286 => x"f8518480",
   287 => x"8082872d",
   288 => x"80578c16",
   289 => x"085574fa",
   290 => x"d5abfddc",
   291 => x"2e93388c",
   292 => x"16085284",
   293 => x"80809cb4",
   294 => x"51848080",
   295 => x"82872d80",
   296 => x"57755580",
   297 => x"74258e38",
   298 => x"74708405",
   299 => x"5608ff15",
   300 => x"555373f4",
   301 => x"38750854",
   302 => x"73fce0c9",
   303 => x"aad52e92",
   304 => x"38750852",
   305 => x"8480809c",
   306 => x"f0518480",
   307 => x"8082872d",
   308 => x"80578c16",
   309 => x"085372fa",
   310 => x"d5abfddc",
   311 => x"2e93388c",
   312 => x"16085284",
   313 => x"80809dac",
   314 => x"51848080",
   315 => x"82872d80",
   316 => x"578f0b82",
   317 => x"1734f00b",
   318 => x"8d173475",
   319 => x"337081ff",
   320 => x"06565474",
   321 => x"81cc2e97",
   322 => x"38753370",
   323 => x"81ff0653",
   324 => x"57848080",
   325 => x"9de85184",
   326 => x"80808287",
   327 => x"2d805781",
   328 => x"16337081",
   329 => x"ff065455",
   330 => x"72922e98",
   331 => x"38811633",
   332 => x"7081ff06",
   333 => x"53548480",
   334 => x"809e9051",
   335 => x"84808082",
   336 => x"872d8057",
   337 => x"82163370",
   338 => x"81ff0654",
   339 => x"55728f2e",
   340 => x"98388216",
   341 => x"337081ff",
   342 => x"06535784",
   343 => x"80809eb8",
   344 => x"51848080",
   345 => x"82872d80",
   346 => x"57831633",
   347 => x"7081ff06",
   348 => x"55537380",
   349 => x"d52e9838",
   350 => x"83163370",
   351 => x"81ff0653",
   352 => x"55848080",
   353 => x"9ee05184",
   354 => x"80808287",
   355 => x"2d80578c",
   356 => x"16337081",
   357 => x"ff065553",
   358 => x"7381aa2e",
   359 => x"98388c16",
   360 => x"337081ff",
   361 => x"06535784",
   362 => x"80809f88",
   363 => x"51848080",
   364 => x"82872d80",
   365 => x"578d1633",
   366 => x"7081ff06",
   367 => x"56547481",
   368 => x"f02e9838",
   369 => x"8d163370",
   370 => x"81ff0653",
   371 => x"53848080",
   372 => x"9fb45184",
   373 => x"80808287",
   374 => x"2d80578e",
   375 => x"16337081",
   376 => x"ff065654",
   377 => x"7481fe2e",
   378 => x"98388e16",
   379 => x"337081ff",
   380 => x"06535784",
   381 => x"80809fe0",
   382 => x"51848080",
   383 => x"82872d80",
   384 => x"578f1633",
   385 => x"7081ff06",
   386 => x"54557281",
   387 => x"dc2e9838",
   388 => x"8f163370",
   389 => x"81ff0653",
   390 => x"54848080",
   391 => x"a08c5184",
   392 => x"80808287",
   393 => x"2d805775",
   394 => x"227083ff",
   395 => x"ff065455",
   396 => x"72839892",
   397 => x"2e983875",
   398 => x"227083ff",
   399 => x"ff065357",
   400 => x"848080a0",
   401 => x"b8518480",
   402 => x"8082872d",
   403 => x"80578e16",
   404 => x"227083ff",
   405 => x"ff065553",
   406 => x"7383fddc",
   407 => x"2e99388e",
   408 => x"16227083",
   409 => x"ffff0653",
   410 => x"55848080",
   411 => x"a0e05184",
   412 => x"80808287",
   413 => x"2d805776",
   414 => x"848080a8",
   415 => x"c40c029c",
   416 => x"050d0402",
   417 => x"e8050d77",
   418 => x"79555680",
   419 => x"c4c4b376",
   420 => x"0c84a2d5",
   421 => x"ccf70b84",
   422 => x"170cf8c4",
   423 => x"e6d5bb0b",
   424 => x"88170cfc",
   425 => x"e6f7ddff",
   426 => x"0b8c170c",
   427 => x"85aad6d5",
   428 => x"aa0b9017",
   429 => x"0c821608",
   430 => x"53728291",
   431 => x"cd88d52e",
   432 => x"8f387252",
   433 => x"848080a1",
   434 => x"88518480",
   435 => x"8082872d",
   436 => x"86160853",
   437 => x"7286b3de",
   438 => x"91992e8f",
   439 => x"38725284",
   440 => x"8080a1c4",
   441 => x"51848080",
   442 => x"82872d8a",
   443 => x"16085372",
   444 => x"fad5ef99",
   445 => x"dd2e8f38",
   446 => x"72528480",
   447 => x"80a28051",
   448 => x"84808082",
   449 => x"872d8e16",
   450 => x"085372fe",
   451 => x"f7fdaad5",
   452 => x"2e8f3872",
   453 => x"52848080",
   454 => x"a2bc5184",
   455 => x"80808287",
   456 => x"2d755580",
   457 => x"74258e38",
   458 => x"74708405",
   459 => x"5608ff15",
   460 => x"555373f4",
   461 => x"38821608",
   462 => x"53728291",
   463 => x"cd88d52e",
   464 => x"8f387252",
   465 => x"848080a2",
   466 => x"f8518480",
   467 => x"8082872d",
   468 => x"86160853",
   469 => x"7286b3de",
   470 => x"91992e8f",
   471 => x"38725284",
   472 => x"8080a3b4",
   473 => x"51848080",
   474 => x"82872d8a",
   475 => x"16085372",
   476 => x"fad5ef99",
   477 => x"dd2e8f38",
   478 => x"72528480",
   479 => x"80a3f051",
   480 => x"84808082",
   481 => x"872d8e16",
   482 => x"085372fe",
   483 => x"f7fdaad5",
   484 => x"2e8f3872",
   485 => x"52848080",
   486 => x"a4ac5184",
   487 => x"80808287",
   488 => x"2d728480",
   489 => x"80a8c40c",
   490 => x"0298050d",
   491 => x"0402cc05",
   492 => x"0d7e5a80",
   493 => x"0b848080",
   494 => x"a4e85259",
   495 => x"84808082",
   496 => x"872d80e1",
   497 => x"b35780fe",
   498 => x"5dae5184",
   499 => x"808085db",
   500 => x"2d765c8f",
   501 => x"ffff5876",
   502 => x"bfffff06",
   503 => x"7010101b",
   504 => x"56750c76",
   505 => x"1070962a",
   506 => x"81065657",
   507 => x"74802e85",
   508 => x"38768107",
   509 => x"5776952a",
   510 => x"81065574",
   511 => x"802e8538",
   512 => x"76813257",
   513 => x"ff185877",
   514 => x"8025cc38",
   515 => x"7b578fff",
   516 => x"ff5876bf",
   517 => x"ffff0670",
   518 => x"10101b70",
   519 => x"08575d56",
   520 => x"74762e81",
   521 => x"8b388079",
   522 => x"53848080",
   523 => x"a4f8525b",
   524 => x"84808082",
   525 => x"872d7454",
   526 => x"75537552",
   527 => x"848080a5",
   528 => x"8c518480",
   529 => x"8082872d",
   530 => x"7a597610",
   531 => x"70962a81",
   532 => x"06565774",
   533 => x"802e8538",
   534 => x"76810757",
   535 => x"76952a81",
   536 => x"065c7b80",
   537 => x"2e853876",
   538 => x"813257ff",
   539 => x"18587780",
   540 => x"25ff9f38",
   541 => x"76107096",
   542 => x"2a810659",
   543 => x"5777802e",
   544 => x"85387681",
   545 => x"07577695",
   546 => x"2a81065c",
   547 => x"7b802e85",
   548 => x"38768132",
   549 => x"57ff1d5d",
   550 => x"7cfeae38",
   551 => x"8a518480",
   552 => x"8085db2d",
   553 => x"7a848080",
   554 => x"a8c40c02",
   555 => x"b4050d04",
   556 => x"81195984",
   557 => x"808090ca",
   558 => x"0402c805",
   559 => x"0d7f5d80",
   560 => x"61922bff",
   561 => x"055b5b80",
   562 => x"e1b30b84",
   563 => x"8080a5b4",
   564 => x"52578480",
   565 => x"8082872d",
   566 => x"7a7a2781",
   567 => x"9e387c7a",
   568 => x"5a587678",
   569 => x"0c761070",
   570 => x"962a7081",
   571 => x"06515757",
   572 => x"75802e85",
   573 => x"38768107",
   574 => x"5776952a",
   575 => x"70810651",
   576 => x"5675802e",
   577 => x"85387681",
   578 => x"3257ff19",
   579 => x"84195959",
   580 => x"78d03880",
   581 => x"e1b35780",
   582 => x"7a2780df",
   583 => x"387c5877",
   584 => x"08567577",
   585 => x"2e80e838",
   586 => x"807b5384",
   587 => x"8080a4f8",
   588 => x"525c8480",
   589 => x"8082872d",
   590 => x"7d557554",
   591 => x"76537852",
   592 => x"848080a5",
   593 => x"c8518480",
   594 => x"8082872d",
   595 => x"7b5b7610",
   596 => x"70962a81",
   597 => x"065e577c",
   598 => x"802e8538",
   599 => x"76810757",
   600 => x"76952a81",
   601 => x"065d7c80",
   602 => x"2e853876",
   603 => x"81325781",
   604 => x"19841959",
   605 => x"59797926",
   606 => x"ffa5388a",
   607 => x"51848080",
   608 => x"85db2d7b",
   609 => x"848080a8",
   610 => x"c40c02b8",
   611 => x"050d0481",
   612 => x"1b5b8480",
   613 => x"8092ce04",
   614 => x"02cc050d",
   615 => x"7e605e58",
   616 => x"815a805b",
   617 => x"80c07a58",
   618 => x"5c85ada9",
   619 => x"89bb780c",
   620 => x"79598156",
   621 => x"97557676",
   622 => x"07822b78",
   623 => x"11515485",
   624 => x"ada989bb",
   625 => x"740c7510",
   626 => x"ff165656",
   627 => x"748025e6",
   628 => x"38761081",
   629 => x"1a5a5798",
   630 => x"7925d738",
   631 => x"7756807d",
   632 => x"2590387c",
   633 => x"55757084",
   634 => x"055708ff",
   635 => x"16565474",
   636 => x"f4388157",
   637 => x"ff8787a5",
   638 => x"c3780c97",
   639 => x"5976822b",
   640 => x"78117008",
   641 => x"5f56567c",
   642 => x"ff8787a5",
   643 => x"c32e80cc",
   644 => x"38740854",
   645 => x"7385ada9",
   646 => x"89bb2e94",
   647 => x"38807508",
   648 => x"54765384",
   649 => x"8080a5fc",
   650 => x"525a8480",
   651 => x"8082872d",
   652 => x"7610ff1a",
   653 => x"5a577880",
   654 => x"25c3387a",
   655 => x"822b5675",
   656 => x"b1387b52",
   657 => x"848080a6",
   658 => x"9c518480",
   659 => x"8082872d",
   660 => x"7b848080",
   661 => x"a8c40c02",
   662 => x"b4050d04",
   663 => x"7a770777",
   664 => x"10ff1b5b",
   665 => x"585b7880",
   666 => x"25ff9238",
   667 => x"84808094",
   668 => x"bb047552",
   669 => x"848080a6",
   670 => x"d8518480",
   671 => x"8082872d",
   672 => x"75992a81",
   673 => x"32810670",
   674 => x"09810571",
   675 => x"07700970",
   676 => x"9f2c7d06",
   677 => x"79109fff",
   678 => x"fffc0660",
   679 => x"812a415a",
   680 => x"5d575859",
   681 => x"75da3879",
   682 => x"09810570",
   683 => x"7b079f2a",
   684 => x"55567bbf",
   685 => x"26843873",
   686 => x"9d388170",
   687 => x"53848080",
   688 => x"a69c525c",
   689 => x"84808082",
   690 => x"872d7b84",
   691 => x"8080a8c4",
   692 => x"0c02b405",
   693 => x"0d048480",
   694 => x"80a6f051",
   695 => x"84808082",
   696 => x"872d7b52",
   697 => x"848080a6",
   698 => x"9c518480",
   699 => x"8082872d",
   700 => x"7b848080",
   701 => x"a8c40c02",
   702 => x"b4050d04",
   703 => x"02cc050d",
   704 => x"810b8480",
   705 => x"8099f05a",
   706 => x"5a835b78",
   707 => x"08800c80",
   708 => x"08790858",
   709 => x"5675772e",
   710 => x"94388008",
   711 => x"53765284",
   712 => x"80809a80",
   713 => x"51848080",
   714 => x"82872d80",
   715 => x"5a807059",
   716 => x"57777084",
   717 => x"05590881",
   718 => x"185856a0",
   719 => x"807724f1",
   720 => x"38800879",
   721 => x"08585877",
   722 => x"772e9438",
   723 => x"80085376",
   724 => x"52848080",
   725 => x"9ac05184",
   726 => x"80808287",
   727 => x"2d805aff",
   728 => x"1b841a5a",
   729 => x"5b7a8025",
   730 => x"ffa13879",
   731 => x"802e8d38",
   732 => x"848080a7",
   733 => x"bc518480",
   734 => x"8082872d",
   735 => x"a0805280",
   736 => x"51848080",
   737 => x"87ed2d84",
   738 => x"8080a8c4",
   739 => x"08802e8d",
   740 => x"38848080",
   741 => x"a7e05184",
   742 => x"80808287",
   743 => x"2da08052",
   744 => x"80518480",
   745 => x"8093982d",
   746 => x"848080a8",
   747 => x"c4085a84",
   748 => x"8080a8c4",
   749 => x"08802e8d",
   750 => x"38848080",
   751 => x"a7fc5184",
   752 => x"80808287",
   753 => x"2d807a90",
   754 => x"808029ff",
   755 => x"055a5b80",
   756 => x"e1b30b84",
   757 => x"8080a5b4",
   758 => x"52578480",
   759 => x"8082872d",
   760 => x"7a587a79",
   761 => x"2781a238",
   762 => x"77822b77",
   763 => x"710c5676",
   764 => x"1070962a",
   765 => x"70810651",
   766 => x"57577580",
   767 => x"2e853876",
   768 => x"81075776",
   769 => x"952a7081",
   770 => x"06515675",
   771 => x"802e8538",
   772 => x"76813257",
   773 => x"81185878",
   774 => x"7826cd38",
   775 => x"80e1b357",
   776 => x"80587779",
   777 => x"2780e238",
   778 => x"77822b70",
   779 => x"08515675",
   780 => x"772e81a0",
   781 => x"38807b53",
   782 => x"848080a4",
   783 => x"f8525c84",
   784 => x"80808287",
   785 => x"2d7c5575",
   786 => x"54765377",
   787 => x"52848080",
   788 => x"a5c85184",
   789 => x"80808287",
   790 => x"2d7b5b76",
   791 => x"1070962a",
   792 => x"70810651",
   793 => x"57577580",
   794 => x"2e853876",
   795 => x"81075776",
   796 => x"952a7081",
   797 => x"06515675",
   798 => x"802e8538",
   799 => x"76813257",
   800 => x"81185878",
   801 => x"7826ffa0",
   802 => x"388a5184",
   803 => x"808085db",
   804 => x"2d7b802e",
   805 => x"8d388480",
   806 => x"80a89451",
   807 => x"84808082",
   808 => x"872d7952",
   809 => x"80518480",
   810 => x"808fad2d",
   811 => x"848080a8",
   812 => x"c408802e",
   813 => x"fcca3884",
   814 => x"8080a8ac",
   815 => x"51848080",
   816 => x"82872d81",
   817 => x"0b848080",
   818 => x"99f05a5a",
   819 => x"835b8480",
   820 => x"80968b04",
   821 => x"811b5b84",
   822 => x"808098db",
   823 => x"04000000",
   824 => x"00ffffff",
   825 => x"ff00ffff",
   826 => x"ffff00ff",
   827 => x"ffffff00",
   828 => x"00000000",
   829 => x"55555555",
   830 => x"aaaaaaaa",
   831 => x"ffffffff",
   832 => x"53616e69",
   833 => x"74792063",
   834 => x"6865636b",
   835 => x"20666169",
   836 => x"6c656420",
   837 => x"28626566",
   838 => x"6f726520",
   839 => x"63616368",
   840 => x"65207265",
   841 => x"66726573",
   842 => x"6829206f",
   843 => x"6e203078",
   844 => x"25642028",
   845 => x"676f7420",
   846 => x"30782564",
   847 => x"290a0000",
   848 => x"53616e69",
   849 => x"74792063",
   850 => x"6865636b",
   851 => x"20666169",
   852 => x"6c656420",
   853 => x"28616674",
   854 => x"65722063",
   855 => x"61636865",
   856 => x"20726566",
   857 => x"72657368",
   858 => x"29206f6e",
   859 => x"20307825",
   860 => x"64202867",
   861 => x"6f742030",
   862 => x"78256429",
   863 => x"0a000000",
   864 => x"42797465",
   865 => x"20636865",
   866 => x"636b2066",
   867 => x"61696c65",
   868 => x"64202862",
   869 => x"65666f72",
   870 => x"65206361",
   871 => x"63686520",
   872 => x"72656672",
   873 => x"65736829",
   874 => x"20617420",
   875 => x"30202867",
   876 => x"6f742030",
   877 => x"78256429",
   878 => x"0a000000",
   879 => x"42797465",
   880 => x"20636865",
   881 => x"636b2066",
   882 => x"61696c65",
   883 => x"64202862",
   884 => x"65666f72",
   885 => x"65206361",
   886 => x"63686520",
   887 => x"72656672",
   888 => x"65736829",
   889 => x"20617420",
   890 => x"33202867",
   891 => x"6f742030",
   892 => x"78256429",
   893 => x"0a000000",
   894 => x"42797465",
   895 => x"20636865",
   896 => x"636b2032",
   897 => x"20666169",
   898 => x"6c656420",
   899 => x"28626566",
   900 => x"6f726520",
   901 => x"63616368",
   902 => x"65207265",
   903 => x"66726573",
   904 => x"68292061",
   905 => x"74203020",
   906 => x"28676f74",
   907 => x"20307825",
   908 => x"64290a00",
   909 => x"42797465",
   910 => x"20636865",
   911 => x"636b2032",
   912 => x"20666169",
   913 => x"6c656420",
   914 => x"28626566",
   915 => x"6f726520",
   916 => x"63616368",
   917 => x"65207265",
   918 => x"66726573",
   919 => x"68292061",
   920 => x"74203320",
   921 => x"28676f74",
   922 => x"20307825",
   923 => x"64290a00",
   924 => x"42797465",
   925 => x"20636865",
   926 => x"636b2066",
   927 => x"61696c65",
   928 => x"64202861",
   929 => x"66746572",
   930 => x"20636163",
   931 => x"68652072",
   932 => x"65667265",
   933 => x"73682920",
   934 => x"61742030",
   935 => x"2028676f",
   936 => x"74203078",
   937 => x"2564290a",
   938 => x"00000000",
   939 => x"42797465",
   940 => x"20636865",
   941 => x"636b2066",
   942 => x"61696c65",
   943 => x"64202861",
   944 => x"66746572",
   945 => x"20636163",
   946 => x"68652072",
   947 => x"65667265",
   948 => x"73682920",
   949 => x"61742033",
   950 => x"2028676f",
   951 => x"74203078",
   952 => x"2564290a",
   953 => x"00000000",
   954 => x"42797465",
   955 => x"20726561",
   956 => x"64206368",
   957 => x"65636b20",
   958 => x"6661696c",
   959 => x"65642061",
   960 => x"74203020",
   961 => x"28676f74",
   962 => x"20307825",
   963 => x"64290a00",
   964 => x"42797465",
   965 => x"20726561",
   966 => x"64206368",
   967 => x"65636b20",
   968 => x"6661696c",
   969 => x"65642061",
   970 => x"74203120",
   971 => x"28676f74",
   972 => x"20307825",
   973 => x"64290a00",
   974 => x"42797465",
   975 => x"20726561",
   976 => x"64206368",
   977 => x"65636b20",
   978 => x"6661696c",
   979 => x"65642061",
   980 => x"74203220",
   981 => x"28676f74",
   982 => x"20307825",
   983 => x"64290a00",
   984 => x"42797465",
   985 => x"20726561",
   986 => x"64206368",
   987 => x"65636b20",
   988 => x"6661696c",
   989 => x"65642061",
   990 => x"74203320",
   991 => x"28676f74",
   992 => x"20307825",
   993 => x"64290a00",
   994 => x"42797465",
   995 => x"20726561",
   996 => x"64206368",
   997 => x"65636b20",
   998 => x"6661696c",
   999 => x"65642061",
  1000 => x"74203132",
  1001 => x"2028676f",
  1002 => x"74203078",
  1003 => x"2564290a",
  1004 => x"00000000",
  1005 => x"42797465",
  1006 => x"20726561",
  1007 => x"64206368",
  1008 => x"65636b20",
  1009 => x"6661696c",
  1010 => x"65642061",
  1011 => x"74203133",
  1012 => x"2028676f",
  1013 => x"74203078",
  1014 => x"2564290a",
  1015 => x"00000000",
  1016 => x"42797465",
  1017 => x"20726561",
  1018 => x"64206368",
  1019 => x"65636b20",
  1020 => x"6661696c",
  1021 => x"65642061",
  1022 => x"74203134",
  1023 => x"2028676f",
  1024 => x"74203078",
  1025 => x"2564290a",
  1026 => x"00000000",
  1027 => x"42797465",
  1028 => x"20726561",
  1029 => x"64206368",
  1030 => x"65636b20",
  1031 => x"6661696c",
  1032 => x"65642061",
  1033 => x"74203135",
  1034 => x"2028676f",
  1035 => x"74203078",
  1036 => x"2564290a",
  1037 => x"00000000",
  1038 => x"576f7264",
  1039 => x"20726561",
  1040 => x"64206368",
  1041 => x"65636b20",
  1042 => x"6661696c",
  1043 => x"65642061",
  1044 => x"74203020",
  1045 => x"28676f74",
  1046 => x"20307825",
  1047 => x"64290a00",
  1048 => x"576f7264",
  1049 => x"20726561",
  1050 => x"64206368",
  1051 => x"65636b20",
  1052 => x"6661696c",
  1053 => x"65642061",
  1054 => x"74203720",
  1055 => x"28676f74",
  1056 => x"20307825",
  1057 => x"64290a00",
  1058 => x"416c6967",
  1059 => x"6e206368",
  1060 => x"65636b20",
  1061 => x"6661696c",
  1062 => x"65642028",
  1063 => x"6265666f",
  1064 => x"72652063",
  1065 => x"61636865",
  1066 => x"20726566",
  1067 => x"72657368",
  1068 => x"29206174",
  1069 => x"20322028",
  1070 => x"676f7420",
  1071 => x"30782564",
  1072 => x"290a0000",
  1073 => x"416c6967",
  1074 => x"6e206368",
  1075 => x"65636b20",
  1076 => x"6661696c",
  1077 => x"65642028",
  1078 => x"6265666f",
  1079 => x"72652063",
  1080 => x"61636865",
  1081 => x"20726566",
  1082 => x"72657368",
  1083 => x"29206174",
  1084 => x"20362028",
  1085 => x"676f7420",
  1086 => x"30782564",
  1087 => x"290a0000",
  1088 => x"416c6967",
  1089 => x"6e206368",
  1090 => x"65636b20",
  1091 => x"6661696c",
  1092 => x"65642028",
  1093 => x"6265666f",
  1094 => x"72652063",
  1095 => x"61636865",
  1096 => x"20726566",
  1097 => x"72657368",
  1098 => x"29206174",
  1099 => x"20313020",
  1100 => x"28676f74",
  1101 => x"20307825",
  1102 => x"64290a00",
  1103 => x"416c6967",
  1104 => x"6e206368",
  1105 => x"65636b20",
  1106 => x"6661696c",
  1107 => x"65642028",
  1108 => x"6265666f",
  1109 => x"72652063",
  1110 => x"61636865",
  1111 => x"20726566",
  1112 => x"72657368",
  1113 => x"29206174",
  1114 => x"20313420",
  1115 => x"28676f74",
  1116 => x"20307825",
  1117 => x"64290a00",
  1118 => x"416c6967",
  1119 => x"6e206368",
  1120 => x"65636b20",
  1121 => x"6661696c",
  1122 => x"65642028",
  1123 => x"61667465",
  1124 => x"72206361",
  1125 => x"63686520",
  1126 => x"72656672",
  1127 => x"65736829",
  1128 => x"20617420",
  1129 => x"32202867",
  1130 => x"6f742030",
  1131 => x"78256429",
  1132 => x"0a000000",
  1133 => x"416c6967",
  1134 => x"6e206368",
  1135 => x"65636b20",
  1136 => x"6661696c",
  1137 => x"65642028",
  1138 => x"61667465",
  1139 => x"72206361",
  1140 => x"63686520",
  1141 => x"72656672",
  1142 => x"65736829",
  1143 => x"20617420",
  1144 => x"36202867",
  1145 => x"6f742030",
  1146 => x"78256429",
  1147 => x"0a000000",
  1148 => x"416c6967",
  1149 => x"6e206368",
  1150 => x"65636b20",
  1151 => x"6661696c",
  1152 => x"65642028",
  1153 => x"61667465",
  1154 => x"72206361",
  1155 => x"63686520",
  1156 => x"72656672",
  1157 => x"65736829",
  1158 => x"20617420",
  1159 => x"31302028",
  1160 => x"676f7420",
  1161 => x"30782564",
  1162 => x"290a0000",
  1163 => x"416c6967",
  1164 => x"6e206368",
  1165 => x"65636b20",
  1166 => x"6661696c",
  1167 => x"65642028",
  1168 => x"61667465",
  1169 => x"72206361",
  1170 => x"63686520",
  1171 => x"72656672",
  1172 => x"65736829",
  1173 => x"20617420",
  1174 => x"31342028",
  1175 => x"676f7420",
  1176 => x"30782564",
  1177 => x"290a0000",
  1178 => x"43686563",
  1179 => x"6b696e67",
  1180 => x"206d656d",
  1181 => x"6f727900",
  1182 => x"30782564",
  1183 => x"20676f6f",
  1184 => x"64207265",
  1185 => x"6164732c",
  1186 => x"20000000",
  1187 => x"4572726f",
  1188 => x"72206174",
  1189 => x"20307825",
  1190 => x"642c2065",
  1191 => x"78706563",
  1192 => x"74656420",
  1193 => x"30782564",
  1194 => x"2c20676f",
  1195 => x"74203078",
  1196 => x"25640a00",
  1197 => x"4c696e65",
  1198 => x"6172206d",
  1199 => x"656d6f72",
  1200 => x"79206368",
  1201 => x"65636b00",
  1202 => x"4572726f",
  1203 => x"72206174",
  1204 => x"20307825",
  1205 => x"642c2065",
  1206 => x"78706563",
  1207 => x"74656420",
  1208 => x"30782564",
  1209 => x"2c20676f",
  1210 => x"74203078",
  1211 => x"2564206f",
  1212 => x"6e20726f",
  1213 => x"756e6420",
  1214 => x"25640a00",
  1215 => x"42616420",
  1216 => x"64617461",
  1217 => x"20666f75",
  1218 => x"6e642061",
  1219 => x"74203078",
  1220 => x"25642028",
  1221 => x"30782564",
  1222 => x"290a0000",
  1223 => x"53445241",
  1224 => x"4d207369",
  1225 => x"7a652028",
  1226 => x"61737375",
  1227 => x"6d696e67",
  1228 => x"206e6f20",
  1229 => x"61646472",
  1230 => x"65737320",
  1231 => x"6661756c",
  1232 => x"74732920",
  1233 => x"69732030",
  1234 => x"78256420",
  1235 => x"6d656761",
  1236 => x"62797465",
  1237 => x"730a0000",
  1238 => x"416c6961",
  1239 => x"73657320",
  1240 => x"666f756e",
  1241 => x"64206174",
  1242 => x"20307825",
  1243 => x"640a0000",
  1244 => x"28416c69",
  1245 => x"61736573",
  1246 => x"2070726f",
  1247 => x"6261626c",
  1248 => x"79207369",
  1249 => x"6d706c79",
  1250 => x"20696e64",
  1251 => x"69636174",
  1252 => x"65207468",
  1253 => x"61742052",
  1254 => x"414d0a69",
  1255 => x"7320736d",
  1256 => x"616c6c65",
  1257 => x"72207468",
  1258 => x"616e2036",
  1259 => x"34206d65",
  1260 => x"67616279",
  1261 => x"74657329",
  1262 => x"0a000000",
  1263 => x"46697273",
  1264 => x"74207374",
  1265 => x"61676520",
  1266 => x"73616e69",
  1267 => x"74792063",
  1268 => x"6865636b",
  1269 => x"20706173",
  1270 => x"7365642e",
  1271 => x"0a000000",
  1272 => x"42797465",
  1273 => x"20286471",
  1274 => x"6d292063",
  1275 => x"6865636b",
  1276 => x"20706173",
  1277 => x"7365640a",
  1278 => x"00000000",
  1279 => x"41646472",
  1280 => x"65737320",
  1281 => x"63686563",
  1282 => x"6b207061",
  1283 => x"73736564",
  1284 => x"2e0a0000",
  1285 => x"4c696e65",
  1286 => x"61722063",
  1287 => x"6865636b",
  1288 => x"20706173",
  1289 => x"7365642e",
  1290 => x"0a0a0000",
  1291 => x"4c465352",
  1292 => x"20636865",
  1293 => x"636b2070",
  1294 => x"61737365",
  1295 => x"642e0a0a",
  1296 => x"00000000",
	others => x"00000000"
);

begin

process (clk)
begin
	if (clk'event and clk = '1') then
		if (from_zpu.memAWriteEnable = '1') and (from_zpu.memBWriteEnable = '1') and (from_zpu.memAAddr=from_zpu.memBAddr) and (from_zpu.memAWrite/=from_zpu.memBWrite) then
			report "write collision" severity failure;
		end if;
	
		if (from_zpu.memAWriteEnable = '1') then
			ram(to_integer(unsigned(from_zpu.memAAddr(maxAddrBitBRAM downto 2)))) := from_zpu.memAWrite;
			to_zpu.memARead <= from_zpu.memAWrite;
		else
			to_zpu.memARead <= ram(to_integer(unsigned(from_zpu.memAAddr(maxAddrBitBRAM downto 2))));
		end if;
	end if;
end process;

process (clk)
begin
	if (clk'event and clk = '1') then
		if (from_zpu.memBWriteEnable = '1') then
			ram(to_integer(unsigned(from_zpu.memBAddr(maxAddrBitBRAM downto 2)))) := from_zpu.memBWrite;
			to_zpu.memBRead <= from_zpu.memBWrite;
		else
			to_zpu.memBRead <= ram(to_integer(unsigned(from_zpu.memBAddr(maxAddrBitBRAM downto 2))));
		end if;
	end if;
end process;


end arch;

