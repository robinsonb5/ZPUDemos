-- ZPU
--
-- Copyright 2004-2008 oharboe - �yvind Harboe - oyvind.harboe@zylin.com
-- Modified by Alastair M. Robinson for the ZPUFlex project.
--
-- The FreeBSD license
-- 
-- Redistribution and use in source and binary forms, with or without
-- modification, are permitted provided that the following conditions
-- are met:
-- 
-- 1. Redistributions of source code must retain the above copyright
--    notice, this list of conditions and the following disclaimer.
-- 2. Redistributions in binary form must reproduce the above
--    copyright notice, this list of conditions and the following
--    disclaimer in the documentation and/or other materials
--    provided with the distribution.
-- 
-- THIS SOFTWARE IS PROVIDED BY THE ZPU PROJECT ``AS IS'' AND ANY
-- EXPRESS OR IMPLIED WARRANTIES, INCLUDING, BUT NOT LIMITED TO,
-- THE IMPLIED WARRANTIES OF MERCHANTABILITY AND FITNESS FOR A
-- PARTICULAR PURPOSE ARE DISCLAIMED. IN NO EVENT SHALL THE
-- ZPU PROJECT OR CONTRIBUTORS BE LIABLE FOR ANY DIRECT,
-- INDIRECT, INCIDENTAL, SPECIAL, EXEMPLARY, OR CONSEQUENTIAL DAMAGES
-- (INCLUDING, BUT NOT LIMITED TO, PROCUREMENT OF SUBSTITUTE GOODS
-- OR SERVICES; LOSS OF USE, DATA, OR PROFITS; OR BUSINESS INTERRUPTION)
-- HOWEVER CAUSED AND ON ANY THEORY OF LIABILITY, WHETHER IN CONTRACT,
-- STRICT LIABILITY, OR TORT (INCLUDING NEGLIGENCE OR OTHERWISE)
-- ARISING IN ANY WAY OUT OF THE USE OF THIS SOFTWARE, EVEN IF
-- ADVISED OF THE POSSIBILITY OF SUCH DAMAGE.
-- 
-- The views and conclusions contained in the software and documentation
-- are those of the authors and should not be interpreted as representing
-- official policies, either expressed or implied, of the ZPU Project.

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;


library work;
use work.zpu_config.all;
use work.zpupkg.all;

entity SDBootstrap_ROM is
generic
	(
		maxAddrBitBRAM : integer := maxAddrBitBRAMLimit -- Specify your actual ROM size to save LEs and unnecessary block RAM usage.
	);
port (
	clk : in std_logic;
	areset : in std_logic := '0';
	from_zpu : in ZPU_ToROM;
	to_zpu : out ZPU_FromROM
);
end SDBootstrap_ROM;

architecture arch of SDBootstrap_ROM is

type ram_type is array(natural range 0 to ((2**(maxAddrBitBRAM+1))/4)-1) of std_logic_vector(wordSize-1 downto 0);

shared variable ram : ram_type :=
(
     0 => x"84808080",
     1 => x"ed040000",
     2 => x"00000000",
     3 => x"84808080",
     4 => x"880d8004",
     5 => x"84808080",
     6 => x"940471fd",
     7 => x"06087283",
     8 => x"06098105",
     9 => x"8205832b",
    10 => x"2a83ffff",
    11 => x"06520471",
    12 => x"fc060872",
    13 => x"83060981",
    14 => x"05830510",
    15 => x"10102a81",
    16 => x"ff065204",
    17 => x"71fc0608",
    18 => x"848080a0",
    19 => x"cc738306",
    20 => x"10100508",
    21 => x"067381ff",
    22 => x"06738306",
    23 => x"09810583",
    24 => x"05101010",
    25 => x"2b0772fc",
    26 => x"060c5151",
    27 => x"04028405",
    28 => x"84808080",
    29 => x"880c8480",
    30 => x"8080940b",
    31 => x"8480808e",
    32 => x"83040000",
    33 => x"02c4050d",
    34 => x"0280c005",
    35 => x"83ffe0e0",
    36 => x"5b568076",
    37 => x"70840558",
    38 => x"08715e5e",
    39 => x"577c7084",
    40 => x"055e0858",
    41 => x"805b7798",
    42 => x"2a78882b",
    43 => x"59547389",
    44 => x"38765e84",
    45 => x"808083e3",
    46 => x"047b802e",
    47 => x"81fd3880",
    48 => x"5c7380e4",
    49 => x"2ea13873",
    50 => x"80e4268e",
    51 => x"387380e3",
    52 => x"2e819a38",
    53 => x"84808082",
    54 => x"fb047380",
    55 => x"f32e80f5",
    56 => x"38848080",
    57 => x"82fb0475",
    58 => x"84177108",
    59 => x"7e5c5557",
    60 => x"52728025",
    61 => x"8e38ad51",
    62 => x"84808083",
    63 => x"ee2d7209",
    64 => x"81055372",
    65 => x"802ebe38",
    66 => x"8755729c",
    67 => x"2a73842b",
    68 => x"54527180",
    69 => x"2e833881",
    70 => x"59897225",
    71 => x"8a38b712",
    72 => x"52848080",
    73 => x"82aa04b0",
    74 => x"12527880",
    75 => x"2e893871",
    76 => x"51848080",
    77 => x"83ee2dff",
    78 => x"15557480",
    79 => x"25cc3884",
    80 => x"808082cd",
    81 => x"04b05184",
    82 => x"808083ee",
    83 => x"2d805384",
    84 => x"80808394",
    85 => x"04758417",
    86 => x"71087054",
    87 => x"5c575284",
    88 => x"80808492",
    89 => x"2d7b5384",
    90 => x"80808394",
    91 => x"04758417",
    92 => x"71085657",
    93 => x"52848080",
    94 => x"83cb04a5",
    95 => x"51848080",
    96 => x"83ee2d73",
    97 => x"51848080",
    98 => x"83ee2d82",
    99 => x"17578480",
   100 => x"8083d604",
   101 => x"72ff1454",
   102 => x"52807225",
   103 => x"b9387970",
   104 => x"81055b84",
   105 => x"808080af",
   106 => x"2d705254",
   107 => x"84808083",
   108 => x"ee2d8117",
   109 => x"57848080",
   110 => x"83940473",
   111 => x"a52e0981",
   112 => x"06893881",
   113 => x"5c848080",
   114 => x"83d60473",
   115 => x"51848080",
   116 => x"83ee2d81",
   117 => x"1757811b",
   118 => x"5b837b25",
   119 => x"fdc83873",
   120 => x"fdbb387d",
   121 => x"83ffe080",
   122 => x"0c02bc05",
   123 => x"0d0402f8",
   124 => x"050d7352",
   125 => x"c0087088",
   126 => x"2a708106",
   127 => x"51515170",
   128 => x"802ef138",
   129 => x"71c00c71",
   130 => x"83ffe080",
   131 => x"0c028805",
   132 => x"0d0402e8",
   133 => x"050d8078",
   134 => x"57557570",
   135 => x"84055708",
   136 => x"53805472",
   137 => x"982a7388",
   138 => x"2b545271",
   139 => x"802ea238",
   140 => x"c0087088",
   141 => x"2a708106",
   142 => x"51515170",
   143 => x"802ef138",
   144 => x"71c00c81",
   145 => x"15811555",
   146 => x"55837425",
   147 => x"d63871ca",
   148 => x"387483ff",
   149 => x"e0800c02",
   150 => x"98050d04",
   151 => x"02f4050d",
   152 => x"d45281ff",
   153 => x"720c7108",
   154 => x"5381ff72",
   155 => x"0c72882b",
   156 => x"83fe8006",
   157 => x"72087081",
   158 => x"ff065152",
   159 => x"5381ff72",
   160 => x"0c727107",
   161 => x"882b7208",
   162 => x"7081ff06",
   163 => x"51525381",
   164 => x"ff720c72",
   165 => x"7107882b",
   166 => x"72087081",
   167 => x"ff067207",
   168 => x"83ffe080",
   169 => x"0c525302",
   170 => x"8c050d04",
   171 => x"02f4050d",
   172 => x"74767181",
   173 => x"ff06d40c",
   174 => x"535383ff",
   175 => x"f1a00885",
   176 => x"3871892b",
   177 => x"5271982a",
   178 => x"d40c7190",
   179 => x"2a7081ff",
   180 => x"06d40c51",
   181 => x"71882a70",
   182 => x"81ff06d4",
   183 => x"0c517181",
   184 => x"ff06d40c",
   185 => x"72902a70",
   186 => x"81ff06d4",
   187 => x"0c51d408",
   188 => x"7081ff06",
   189 => x"515182b8",
   190 => x"bf527081",
   191 => x"ff2e0981",
   192 => x"06943881",
   193 => x"ff0bd40c",
   194 => x"d4087081",
   195 => x"ff06ff14",
   196 => x"54515171",
   197 => x"e5387083",
   198 => x"ffe0800c",
   199 => x"028c050d",
   200 => x"0402fc05",
   201 => x"0d81c751",
   202 => x"81ff0bd4",
   203 => x"0cff1151",
   204 => x"708025f4",
   205 => x"38028405",
   206 => x"0d0402f0",
   207 => x"050d8480",
   208 => x"8086a12d",
   209 => x"819c9f53",
   210 => x"805287fc",
   211 => x"80f75184",
   212 => x"808085ac",
   213 => x"2d83ffe0",
   214 => x"80085483",
   215 => x"ffe08008",
   216 => x"812e0981",
   217 => x"06ae3881",
   218 => x"ff0bd40c",
   219 => x"820a5284",
   220 => x"9c80e951",
   221 => x"84808085",
   222 => x"ac2d83ff",
   223 => x"e080088e",
   224 => x"3881ff0b",
   225 => x"d40c7353",
   226 => x"84808087",
   227 => x"9b048480",
   228 => x"8086a12d",
   229 => x"ff135372",
   230 => x"ffae3872",
   231 => x"83ffe080",
   232 => x"0c029005",
   233 => x"0d0402f4",
   234 => x"050d81ff",
   235 => x"0bd40c84",
   236 => x"8080a0dc",
   237 => x"51848080",
   238 => x"84922d93",
   239 => x"53805287",
   240 => x"fc80c151",
   241 => x"84808085",
   242 => x"ac2d83ff",
   243 => x"e080088e",
   244 => x"3881ff0b",
   245 => x"d40c8153",
   246 => x"84808087",
   247 => x"ea048480",
   248 => x"8086a12d",
   249 => x"ff135372",
   250 => x"d4387283",
   251 => x"ffe0800c",
   252 => x"028c050d",
   253 => x"0402f005",
   254 => x"0d848080",
   255 => x"86a12d83",
   256 => x"aa52849c",
   257 => x"80c85184",
   258 => x"808085ac",
   259 => x"2d83ffe0",
   260 => x"800883ff",
   261 => x"e0800853",
   262 => x"848080a0",
   263 => x"e8525384",
   264 => x"80808184",
   265 => x"2d72812e",
   266 => x"098106a9",
   267 => x"38848080",
   268 => x"84dc2d83",
   269 => x"ffe08008",
   270 => x"83ffff06",
   271 => x"537283aa",
   272 => x"2ebb3883",
   273 => x"ffe08008",
   274 => x"52848080",
   275 => x"a1805184",
   276 => x"80808184",
   277 => x"2d848080",
   278 => x"87a62d84",
   279 => x"808088f5",
   280 => x"04815484",
   281 => x"80808aa0",
   282 => x"04848080",
   283 => x"a1985184",
   284 => x"80808184",
   285 => x"2d805484",
   286 => x"80808aa0",
   287 => x"0481ff0b",
   288 => x"d40cb153",
   289 => x"84808086",
   290 => x"ba2d83ff",
   291 => x"e0800880",
   292 => x"2e80fe38",
   293 => x"805287fc",
   294 => x"80fa5184",
   295 => x"808085ac",
   296 => x"2d83ffe0",
   297 => x"800880d7",
   298 => x"3883ffe0",
   299 => x"80085284",
   300 => x"8080a1b4",
   301 => x"51848080",
   302 => x"81842d81",
   303 => x"ff0bd40c",
   304 => x"d4087081",
   305 => x"ff067054",
   306 => x"848080a1",
   307 => x"c0535153",
   308 => x"84808081",
   309 => x"842d81ff",
   310 => x"0bd40c81",
   311 => x"ff0bd40c",
   312 => x"81ff0bd4",
   313 => x"0c81ff0b",
   314 => x"d40c7286",
   315 => x"2a708106",
   316 => x"70565153",
   317 => x"72802ea8",
   318 => x"38848080",
   319 => x"88e10483",
   320 => x"ffe08008",
   321 => x"52848080",
   322 => x"a1b45184",
   323 => x"80808184",
   324 => x"2d72822e",
   325 => x"fed338ff",
   326 => x"135372fe",
   327 => x"e7387254",
   328 => x"7383ffe0",
   329 => x"800c0290",
   330 => x"050d0402",
   331 => x"f4050d81",
   332 => x"0b83fff1",
   333 => x"a00cd008",
   334 => x"708f2a70",
   335 => x"81065151",
   336 => x"5372f338",
   337 => x"72d00c84",
   338 => x"808086a1",
   339 => x"2dd00870",
   340 => x"8f2a7081",
   341 => x"06515153",
   342 => x"72f33881",
   343 => x"0bd00c87",
   344 => x"53805284",
   345 => x"d480c051",
   346 => x"84808085",
   347 => x"ac2d83ff",
   348 => x"e0800881",
   349 => x"2e973872",
   350 => x"822e0981",
   351 => x"06893880",
   352 => x"53848080",
   353 => x"8bc704ff",
   354 => x"135372d5",
   355 => x"38848080",
   356 => x"87f52d83",
   357 => x"ffe08008",
   358 => x"83fff1a0",
   359 => x"0c815287",
   360 => x"fc80d051",
   361 => x"84808085",
   362 => x"ac2d81ff",
   363 => x"0bd40cd0",
   364 => x"08708f2a",
   365 => x"70810651",
   366 => x"515372f3",
   367 => x"3872d00c",
   368 => x"81ff0bd4",
   369 => x"0c815372",
   370 => x"83ffe080",
   371 => x"0c028c05",
   372 => x"0d04800b",
   373 => x"83ffe080",
   374 => x"0c0402e0",
   375 => x"050d797b",
   376 => x"57578058",
   377 => x"81ff0bd4",
   378 => x"0cd00870",
   379 => x"8f2a7081",
   380 => x"06515154",
   381 => x"73f33882",
   382 => x"810bd00c",
   383 => x"81ff0bd4",
   384 => x"0c765287",
   385 => x"fc80d151",
   386 => x"84808085",
   387 => x"ac2d80db",
   388 => x"c6df5583",
   389 => x"ffe08008",
   390 => x"802e9b38",
   391 => x"83ffe080",
   392 => x"08537652",
   393 => x"848080a1",
   394 => x"d0518480",
   395 => x"8081842d",
   396 => x"8480808d",
   397 => x"8c0481ff",
   398 => x"0bd40cd4",
   399 => x"087081ff",
   400 => x"06515473",
   401 => x"81fe2e09",
   402 => x"8106a538",
   403 => x"80ff5484",
   404 => x"808084dc",
   405 => x"2d83ffe0",
   406 => x"80087670",
   407 => x"8405580c",
   408 => x"ff145473",
   409 => x"8025e838",
   410 => x"81588480",
   411 => x"808cf604",
   412 => x"ff155574",
   413 => x"c13881ff",
   414 => x"0bd40cd0",
   415 => x"08708f2a",
   416 => x"70810651",
   417 => x"515473f3",
   418 => x"3873d00c",
   419 => x"7783ffe0",
   420 => x"800c02a0",
   421 => x"050d0402",
   422 => x"f4050d74",
   423 => x"70882a83",
   424 => x"fe800670",
   425 => x"72982a07",
   426 => x"72882b87",
   427 => x"fc808006",
   428 => x"73982b81",
   429 => x"f00a0671",
   430 => x"73070783",
   431 => x"ffe0800c",
   432 => x"56515351",
   433 => x"028c050d",
   434 => x"0402f805",
   435 => x"0d028e05",
   436 => x"84808080",
   437 => x"af2d7498",
   438 => x"2b71902b",
   439 => x"0770902c",
   440 => x"83ffe080",
   441 => x"0c525202",
   442 => x"88050d04",
   443 => x"02f8050d",
   444 => x"7370902b",
   445 => x"71902a07",
   446 => x"83ffe080",
   447 => x"0c520288",
   448 => x"050d0402",
   449 => x"ec050d80",
   450 => x"0bfc800c",
   451 => x"848080a1",
   452 => x"f0518480",
   453 => x"8084922d",
   454 => x"8480808a",
   455 => x"ab2d83ff",
   456 => x"e0800880",
   457 => x"2e81f738",
   458 => x"848080a2",
   459 => x"88518480",
   460 => x"8084922d",
   461 => x"84808091",
   462 => x"822d83ff",
   463 => x"e1a05284",
   464 => x"8080a2a0",
   465 => x"51848080",
   466 => x"9de52d83",
   467 => x"ffe08008",
   468 => x"802e81ca",
   469 => x"3883ffe1",
   470 => x"a00b8480",
   471 => x"80a2ac52",
   472 => x"54848080",
   473 => x"84922d80",
   474 => x"55737081",
   475 => x"05558480",
   476 => x"8080af2d",
   477 => x"5372a02e",
   478 => x"80e33872",
   479 => x"a32e8184",
   480 => x"387280c7",
   481 => x"2e098106",
   482 => x"8d388480",
   483 => x"80808c2d",
   484 => x"8480808f",
   485 => x"b804728a",
   486 => x"2e098106",
   487 => x"8d388480",
   488 => x"8080942d",
   489 => x"8480808f",
   490 => x"b8047280",
   491 => x"cc2e0981",
   492 => x"06863883",
   493 => x"ffe1a054",
   494 => x"7281df06",
   495 => x"f0057081",
   496 => x"ff065153",
   497 => x"b8732789",
   498 => x"38ef1370",
   499 => x"81ff0651",
   500 => x"5374842b",
   501 => x"73075584",
   502 => x"80808ee9",
   503 => x"0472a32e",
   504 => x"a3387370",
   505 => x"81055584",
   506 => x"808080af",
   507 => x"2d5372a0",
   508 => x"2ef038ff",
   509 => x"14755370",
   510 => x"52548480",
   511 => x"809de52d",
   512 => x"74fc800c",
   513 => x"73708105",
   514 => x"55848080",
   515 => x"80af2d53",
   516 => x"728a2e09",
   517 => x"8106ed38",
   518 => x"8480808e",
   519 => x"e7048480",
   520 => x"80a2c051",
   521 => x"84808084",
   522 => x"922d800b",
   523 => x"83ffe080",
   524 => x"0c029405",
   525 => x"0d0402e8",
   526 => x"050d7779",
   527 => x"7b585555",
   528 => x"80537276",
   529 => x"25af3874",
   530 => x"70810556",
   531 => x"84808080",
   532 => x"af2d7470",
   533 => x"81055684",
   534 => x"808080af",
   535 => x"2d525271",
   536 => x"712e8938",
   537 => x"81518480",
   538 => x"8090f704",
   539 => x"81135384",
   540 => x"808090c2",
   541 => x"04805170",
   542 => x"83ffe080",
   543 => x"0c029805",
   544 => x"0d0402d8",
   545 => x"050dff0b",
   546 => x"83fff5cc",
   547 => x"0c800b83",
   548 => x"fff5e00c",
   549 => x"848080a2",
   550 => x"cc518480",
   551 => x"8084922d",
   552 => x"83fff1b8",
   553 => x"52805184",
   554 => x"80808bda",
   555 => x"2d83ffe0",
   556 => x"80085483",
   557 => x"ffe08008",
   558 => x"95388480",
   559 => x"80a2dc51",
   560 => x"84808084",
   561 => x"922d7355",
   562 => x"84808099",
   563 => x"a7048480",
   564 => x"80a2f051",
   565 => x"84808084",
   566 => x"922d8056",
   567 => x"810b83ff",
   568 => x"f1ac0c88",
   569 => x"53848080",
   570 => x"a3885283",
   571 => x"fff1ee51",
   572 => x"84808090",
   573 => x"b62d83ff",
   574 => x"e0800876",
   575 => x"2e098106",
   576 => x"8b3883ff",
   577 => x"e0800883",
   578 => x"fff1ac0c",
   579 => x"88538480",
   580 => x"80a39452",
   581 => x"83fff28a",
   582 => x"51848080",
   583 => x"90b62d83",
   584 => x"ffe08008",
   585 => x"8b3883ff",
   586 => x"e0800883",
   587 => x"fff1ac0c",
   588 => x"83fff1ac",
   589 => x"08528480",
   590 => x"80a3a051",
   591 => x"84808081",
   592 => x"842d83ff",
   593 => x"f1ac0880",
   594 => x"2e81cb38",
   595 => x"83fff4fe",
   596 => x"0b848080",
   597 => x"80af2d83",
   598 => x"fff4ff0b",
   599 => x"84808080",
   600 => x"af2d7198",
   601 => x"2b71902b",
   602 => x"0783fff5",
   603 => x"800b8480",
   604 => x"8080af2d",
   605 => x"70882b72",
   606 => x"0783fff5",
   607 => x"810b8480",
   608 => x"8080af2d",
   609 => x"710783ff",
   610 => x"f5b60b84",
   611 => x"808080af",
   612 => x"2d83fff5",
   613 => x"b70b8480",
   614 => x"8080af2d",
   615 => x"71882b07",
   616 => x"535f5452",
   617 => x"5a565755",
   618 => x"7381abaa",
   619 => x"2e098106",
   620 => x"95387551",
   621 => x"8480808d",
   622 => x"972d83ff",
   623 => x"e0800856",
   624 => x"84808093",
   625 => x"df047382",
   626 => x"d4d52e93",
   627 => x"38848080",
   628 => x"a3b45184",
   629 => x"80808492",
   630 => x"2d848080",
   631 => x"95eb0475",
   632 => x"52848080",
   633 => x"a3d45184",
   634 => x"80808184",
   635 => x"2d83fff1",
   636 => x"b8527551",
   637 => x"8480808b",
   638 => x"da2d83ff",
   639 => x"e0800855",
   640 => x"83ffe080",
   641 => x"08802e85",
   642 => x"9e388480",
   643 => x"80a3ec51",
   644 => x"84808084",
   645 => x"922d8480",
   646 => x"80a49451",
   647 => x"84808081",
   648 => x"842d8853",
   649 => x"848080a3",
   650 => x"945283ff",
   651 => x"f28a5184",
   652 => x"808090b6",
   653 => x"2d83ffe0",
   654 => x"80088e38",
   655 => x"810b83ff",
   656 => x"f5e00c84",
   657 => x"808094f7",
   658 => x"04885384",
   659 => x"8080a388",
   660 => x"5283fff1",
   661 => x"ee518480",
   662 => x"8090b62d",
   663 => x"83ffe080",
   664 => x"08802e93",
   665 => x"38848080",
   666 => x"a4ac5184",
   667 => x"80808184",
   668 => x"2d848080",
   669 => x"95eb0483",
   670 => x"fff5b60b",
   671 => x"84808080",
   672 => x"af2d5473",
   673 => x"80d52e09",
   674 => x"810680df",
   675 => x"3883fff5",
   676 => x"b70b8480",
   677 => x"8080af2d",
   678 => x"547381aa",
   679 => x"2e098106",
   680 => x"80c93880",
   681 => x"0b83fff1",
   682 => x"b80b8480",
   683 => x"8080af2d",
   684 => x"56547481",
   685 => x"e92e8338",
   686 => x"81547481",
   687 => x"eb2e8c38",
   688 => x"80557375",
   689 => x"2e098106",
   690 => x"83dd3883",
   691 => x"fff1c30b",
   692 => x"84808080",
   693 => x"af2d5574",
   694 => x"923883ff",
   695 => x"f1c40b84",
   696 => x"808080af",
   697 => x"2d547382",
   698 => x"2e893880",
   699 => x"55848080",
   700 => x"99a70483",
   701 => x"fff1c50b",
   702 => x"84808080",
   703 => x"af2d7083",
   704 => x"fff5e80c",
   705 => x"ff0583ff",
   706 => x"f5dc0c83",
   707 => x"fff1c60b",
   708 => x"84808080",
   709 => x"af2d83ff",
   710 => x"f1c70b84",
   711 => x"808080af",
   712 => x"2d587605",
   713 => x"77828029",
   714 => x"057083ff",
   715 => x"f5d00c83",
   716 => x"fff1c80b",
   717 => x"84808080",
   718 => x"af2d7083",
   719 => x"fff5c80c",
   720 => x"83fff5e0",
   721 => x"08595758",
   722 => x"76802e81",
   723 => x"ea388853",
   724 => x"848080a3",
   725 => x"945283ff",
   726 => x"f28a5184",
   727 => x"808090b6",
   728 => x"2d83ffe0",
   729 => x"800882bf",
   730 => x"3883fff5",
   731 => x"e8087084",
   732 => x"2b83fff5",
   733 => x"b80c7083",
   734 => x"fff5e40c",
   735 => x"83fff1dd",
   736 => x"0b848080",
   737 => x"80af2d83",
   738 => x"fff1dc0b",
   739 => x"84808080",
   740 => x"af2d7182",
   741 => x"80290583",
   742 => x"fff1de0b",
   743 => x"84808080",
   744 => x"af2d7084",
   745 => x"80802912",
   746 => x"83fff1df",
   747 => x"0b848080",
   748 => x"80af2d70",
   749 => x"81800a29",
   750 => x"127083ff",
   751 => x"f1b00c83",
   752 => x"fff5c808",
   753 => x"712983ff",
   754 => x"f5d00805",
   755 => x"7083fff5",
   756 => x"f00c83ff",
   757 => x"f1e50b84",
   758 => x"808080af",
   759 => x"2d83fff1",
   760 => x"e40b8480",
   761 => x"8080af2d",
   762 => x"71828029",
   763 => x"0583fff1",
   764 => x"e60b8480",
   765 => x"8080af2d",
   766 => x"70848080",
   767 => x"291283ff",
   768 => x"f1e70b84",
   769 => x"808080af",
   770 => x"2d70982b",
   771 => x"81f00a06",
   772 => x"72057083",
   773 => x"fff1b40c",
   774 => x"fe117e29",
   775 => x"770583ff",
   776 => x"f5d80c52",
   777 => x"59524354",
   778 => x"5e515259",
   779 => x"525d5759",
   780 => x"57848080",
   781 => x"99a50483",
   782 => x"fff1ca0b",
   783 => x"84808080",
   784 => x"af2d83ff",
   785 => x"f1c90b84",
   786 => x"808080af",
   787 => x"2d718280",
   788 => x"29057083",
   789 => x"fff5b80c",
   790 => x"70a02983",
   791 => x"ff057089",
   792 => x"2a7083ff",
   793 => x"f5e40c83",
   794 => x"fff1cf0b",
   795 => x"84808080",
   796 => x"af2d83ff",
   797 => x"f1ce0b84",
   798 => x"808080af",
   799 => x"2d718280",
   800 => x"29057083",
   801 => x"fff1b00c",
   802 => x"7b71291e",
   803 => x"7083fff5",
   804 => x"d80c7d83",
   805 => x"fff1b40c",
   806 => x"730583ff",
   807 => x"f5f00c55",
   808 => x"5e515155",
   809 => x"55815574",
   810 => x"83ffe080",
   811 => x"0c02a805",
   812 => x"0d0402ec",
   813 => x"050d7670",
   814 => x"872c7180",
   815 => x"ff065755",
   816 => x"5383fff5",
   817 => x"e0088a38",
   818 => x"72882c73",
   819 => x"81ff0656",
   820 => x"547383ff",
   821 => x"f5cc082e",
   822 => x"a93883ff",
   823 => x"f1b85283",
   824 => x"fff5d008",
   825 => x"14518480",
   826 => x"808bda2d",
   827 => x"83ffe080",
   828 => x"085383ff",
   829 => x"e0800880",
   830 => x"2e80cf38",
   831 => x"7383fff5",
   832 => x"cc0c83ff",
   833 => x"f5e00880",
   834 => x"2ea23874",
   835 => x"842983ff",
   836 => x"f1b80570",
   837 => x"08525384",
   838 => x"80808d97",
   839 => x"2d83ffe0",
   840 => x"8008f00a",
   841 => x"06558480",
   842 => x"809ac804",
   843 => x"741083ff",
   844 => x"f1b80570",
   845 => x"84808080",
   846 => x"9a2d5253",
   847 => x"8480808d",
   848 => x"c92d83ff",
   849 => x"e0800855",
   850 => x"74537283",
   851 => x"ffe0800c",
   852 => x"0294050d",
   853 => x"0402cc05",
   854 => x"0d7e605e",
   855 => x"5b8056ff",
   856 => x"0b83fff5",
   857 => x"cc0c83ff",
   858 => x"f1b40883",
   859 => x"fff5d808",
   860 => x"565783ff",
   861 => x"f5e00876",
   862 => x"2e8f3883",
   863 => x"fff5e808",
   864 => x"842b5984",
   865 => x"80809b91",
   866 => x"0483fff5",
   867 => x"e408842b",
   868 => x"59805a79",
   869 => x"792781f0",
   870 => x"38798f06",
   871 => x"a0175754",
   872 => x"73a43874",
   873 => x"52848080",
   874 => x"a4cc5184",
   875 => x"80808184",
   876 => x"2d83fff1",
   877 => x"b8527451",
   878 => x"81155584",
   879 => x"80808bda",
   880 => x"2d83fff1",
   881 => x"b8568076",
   882 => x"84808080",
   883 => x"af2d5558",
   884 => x"73782e83",
   885 => x"38815873",
   886 => x"81e52e81",
   887 => x"a2388170",
   888 => x"7906555c",
   889 => x"73802e81",
   890 => x"96388b16",
   891 => x"84808080",
   892 => x"af2d9806",
   893 => x"58778187",
   894 => x"388b537c",
   895 => x"52755184",
   896 => x"808090b6",
   897 => x"2d83ffe0",
   898 => x"800880f3",
   899 => x"389c1608",
   900 => x"51848080",
   901 => x"8d972d83",
   902 => x"ffe08008",
   903 => x"841c0c9a",
   904 => x"16848080",
   905 => x"809a2d51",
   906 => x"8480808d",
   907 => x"c92d83ff",
   908 => x"e0800883",
   909 => x"ffe08008",
   910 => x"555583ff",
   911 => x"f5e00880",
   912 => x"2ea03894",
   913 => x"16848080",
   914 => x"809a2d51",
   915 => x"8480808d",
   916 => x"c92d83ff",
   917 => x"e0800890",
   918 => x"2b83fff0",
   919 => x"0a067016",
   920 => x"51547388",
   921 => x"1c0c777b",
   922 => x"0c7c5284",
   923 => x"8080a4ec",
   924 => x"51848080",
   925 => x"81842d7b",
   926 => x"54848080",
   927 => x"9dda0481",
   928 => x"1a5a8480",
   929 => x"809b9304",
   930 => x"83fff5e0",
   931 => x"08802e80",
   932 => x"c7387651",
   933 => x"84808099",
   934 => x"b22d83ff",
   935 => x"e0800883",
   936 => x"ffe08008",
   937 => x"53848080",
   938 => x"a5805257",
   939 => x"84808081",
   940 => x"842d7680",
   941 => x"fffffff8",
   942 => x"06547380",
   943 => x"fffffff8",
   944 => x"2e9638fe",
   945 => x"1783fff5",
   946 => x"e8082983",
   947 => x"fff5f008",
   948 => x"05558480",
   949 => x"809b9104",
   950 => x"80547383",
   951 => x"ffe0800c",
   952 => x"02b4050d",
   953 => x"0402e405",
   954 => x"0d787a71",
   955 => x"5483fff5",
   956 => x"bc535555",
   957 => x"8480809a",
   958 => x"d52d83ff",
   959 => x"e0800881",
   960 => x"ff065372",
   961 => x"802e8188",
   962 => x"38848080",
   963 => x"a5985184",
   964 => x"80808492",
   965 => x"2d83fff5",
   966 => x"c00883ff",
   967 => x"05892a57",
   968 => x"80705656",
   969 => x"75772581",
   970 => x"873883ff",
   971 => x"f5c408fe",
   972 => x"0583fff5",
   973 => x"e8082983",
   974 => x"fff5f008",
   975 => x"117683ff",
   976 => x"f5dc0806",
   977 => x"05755452",
   978 => x"53848080",
   979 => x"8bda2d83",
   980 => x"ffe08008",
   981 => x"802e80cc",
   982 => x"38811570",
   983 => x"83fff5dc",
   984 => x"08065455",
   985 => x"72973883",
   986 => x"fff5c408",
   987 => x"51848080",
   988 => x"99b22d83",
   989 => x"ffe08008",
   990 => x"83fff5c4",
   991 => x"0c848014",
   992 => x"81175754",
   993 => x"767624ff",
   994 => x"a1388480",
   995 => x"809fb004",
   996 => x"74528480",
   997 => x"80a5b451",
   998 => x"84808081",
   999 => x"842d8480",
  1000 => x"809fb204",
  1001 => x"83ffe080",
  1002 => x"08538480",
  1003 => x"809fb204",
  1004 => x"81537283",
  1005 => x"ffe0800c",
  1006 => x"029c050d",
  1007 => x"0483ffe0",
  1008 => x"8c080283",
  1009 => x"ffe08c0c",
  1010 => x"ff3d0d80",
  1011 => x"0b83ffe0",
  1012 => x"8c08fc05",
  1013 => x"0c83ffe0",
  1014 => x"8c088805",
  1015 => x"088106ff",
  1016 => x"11700970",
  1017 => x"83ffe08c",
  1018 => x"088c0508",
  1019 => x"0683ffe0",
  1020 => x"8c08fc05",
  1021 => x"081183ff",
  1022 => x"e08c08fc",
  1023 => x"050c83ff",
  1024 => x"e08c0888",
  1025 => x"0508812a",
  1026 => x"83ffe08c",
  1027 => x"0888050c",
  1028 => x"83ffe08c",
  1029 => x"088c0508",
  1030 => x"1083ffe0",
  1031 => x"8c088c05",
  1032 => x"0c515151",
  1033 => x"5183ffe0",
  1034 => x"8c088805",
  1035 => x"08802e84",
  1036 => x"38ffa239",
  1037 => x"83ffe08c",
  1038 => x"08fc0508",
  1039 => x"7083ffe0",
  1040 => x"800c5183",
  1041 => x"3d0d83ff",
  1042 => x"e08c0c04",
  1043 => x"00ffffff",
  1044 => x"ff00ffff",
  1045 => x"ffff00ff",
  1046 => x"ffffff00",
  1047 => x"436d645f",
  1048 => x"696e6974",
  1049 => x"0a000000",
  1050 => x"636d645f",
  1051 => x"434d4438",
  1052 => x"20726573",
  1053 => x"706f6e73",
  1054 => x"653a2025",
  1055 => x"640a0000",
  1056 => x"434d4438",
  1057 => x"5f342072",
  1058 => x"6573706f",
  1059 => x"6e73653a",
  1060 => x"2025640a",
  1061 => x"00000000",
  1062 => x"53444843",
  1063 => x"20496e69",
  1064 => x"7469616c",
  1065 => x"697a6174",
  1066 => x"696f6e20",
  1067 => x"6572726f",
  1068 => x"72210a00",
  1069 => x"434d4435",
  1070 => x"38202564",
  1071 => x"0a202000",
  1072 => x"434d4435",
  1073 => x"385f3220",
  1074 => x"25640a20",
  1075 => x"20000000",
  1076 => x"52656164",
  1077 => x"20636f6d",
  1078 => x"6d616e64",
  1079 => x"20666169",
  1080 => x"6c656420",
  1081 => x"61742025",
  1082 => x"64202825",
  1083 => x"64290a00",
  1084 => x"496e6974",
  1085 => x"69616c69",
  1086 => x"7a696e67",
  1087 => x"20534420",
  1088 => x"63617264",
  1089 => x"0a000000",
  1090 => x"48756e74",
  1091 => x"696e6720",
  1092 => x"666f7220",
  1093 => x"70617274",
  1094 => x"6974696f",
  1095 => x"6e0a0000",
  1096 => x"4d414e49",
  1097 => x"46455354",
  1098 => x"4d535400",
  1099 => x"50617273",
  1100 => x"696e6720",
  1101 => x"6d616e69",
  1102 => x"66657374",
  1103 => x"0a000000",
  1104 => x"52657475",
  1105 => x"726e696e",
  1106 => x"670a0000",
  1107 => x"52656164",
  1108 => x"696e6720",
  1109 => x"4d42520a",
  1110 => x"00000000",
  1111 => x"52656164",
  1112 => x"206f6620",
  1113 => x"4d425220",
  1114 => x"6661696c",
  1115 => x"65640a00",
  1116 => x"4d425220",
  1117 => x"73756363",
  1118 => x"65737366",
  1119 => x"756c6c79",
  1120 => x"20726561",
  1121 => x"640a0000",
  1122 => x"46415431",
  1123 => x"36202020",
  1124 => x"00000000",
  1125 => x"46415433",
  1126 => x"32202020",
  1127 => x"00000000",
  1128 => x"50617274",
  1129 => x"6974696f",
  1130 => x"6e636f75",
  1131 => x"6e742025",
  1132 => x"640a0000",
  1133 => x"4e6f2070",
  1134 => x"61727469",
  1135 => x"74696f6e",
  1136 => x"20736967",
  1137 => x"6e617475",
  1138 => x"72652066",
  1139 => x"6f756e64",
  1140 => x"0a000000",
  1141 => x"52656164",
  1142 => x"696e6720",
  1143 => x"626f6f74",
  1144 => x"20736563",
  1145 => x"746f7220",
  1146 => x"25640a00",
  1147 => x"52656164",
  1148 => x"20626f6f",
  1149 => x"74207365",
  1150 => x"63746f72",
  1151 => x"2066726f",
  1152 => x"6d206669",
  1153 => x"72737420",
  1154 => x"70617274",
  1155 => x"6974696f",
  1156 => x"6e0a0000",
  1157 => x"48756e74",
  1158 => x"696e6720",
  1159 => x"666f7220",
  1160 => x"66696c65",
  1161 => x"73797374",
  1162 => x"656d0a00",
  1163 => x"556e7375",
  1164 => x"70706f72",
  1165 => x"74656420",
  1166 => x"70617274",
  1167 => x"6974696f",
  1168 => x"6e207479",
  1169 => x"7065210d",
  1170 => x"00000000",
  1171 => x"52656164",
  1172 => x"696e6720",
  1173 => x"64697265",
  1174 => x"63746f72",
  1175 => x"79207365",
  1176 => x"63746f72",
  1177 => x"2025640a",
  1178 => x"00000000",
  1179 => x"66696c65",
  1180 => x"20222573",
  1181 => x"2220666f",
  1182 => x"756e640d",
  1183 => x"00000000",
  1184 => x"47657446",
  1185 => x"41544c69",
  1186 => x"6e6b2072",
  1187 => x"65747572",
  1188 => x"6e656420",
  1189 => x"25640a00",
  1190 => x"4f70656e",
  1191 => x"65642066",
  1192 => x"696c652c",
  1193 => x"206c6f61",
  1194 => x"64696e67",
  1195 => x"2e2e2e0a",
  1196 => x"00000000",
  1197 => x"43616e27",
  1198 => x"74206f70",
  1199 => x"656e2025",
  1200 => x"730a0000",
	others => x"00000000"
);

begin

process (clk)
begin
	if (clk'event and clk = '1') then
		if (from_zpu.memAWriteEnable = '1') and (from_zpu.memBWriteEnable = '1') and (from_zpu.memAAddr=from_zpu.memBAddr) and (from_zpu.memAWrite/=from_zpu.memBWrite) then
			report "write collision" severity failure;
		end if;
	
		if (from_zpu.memAWriteEnable = '1') then
			ram(to_integer(unsigned(from_zpu.memAAddr(maxAddrBitBRAM downto 2)))) := from_zpu.memAWrite;
			to_zpu.memARead <= from_zpu.memAWrite;
		else
			to_zpu.memARead <= ram(to_integer(unsigned(from_zpu.memAAddr(maxAddrBitBRAM downto 2))));
		end if;
	end if;
end process;

process (clk)
begin
	if (clk'event and clk = '1') then
		if (from_zpu.memBWriteEnable = '1') then
			ram(to_integer(unsigned(from_zpu.memBAddr(maxAddrBitBRAM downto 2)))) := from_zpu.memBWrite;
			to_zpu.memBRead <= from_zpu.memBWrite;
		else
			to_zpu.memBRead <= ram(to_integer(unsigned(from_zpu.memBAddr(maxAddrBitBRAM downto 2))));
		end if;
	end if;
end process;


end arch;

