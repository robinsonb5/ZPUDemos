-- ZPU
--
-- Copyright 2004-2008 oharboe - �yvind Harboe - oyvind.harboe@zylin.com
-- Modified by Alastair M. Robinson for the ZPUFlex project.
--
-- The FreeBSD license
-- 
-- Redistribution and use in source and binary forms, with or without
-- modification, are permitted provided that the following conditions
-- are met:
-- 
-- 1. Redistributions of source code must retain the above copyright
--    notice, this list of conditions and the following disclaimer.
-- 2. Redistributions in binary form must reproduce the above
--    copyright notice, this list of conditions and the following
--    disclaimer in the documentation and/or other materials
--    provided with the distribution.
-- 
-- THIS SOFTWARE IS PROVIDED BY THE ZPU PROJECT ``AS IS'' AND ANY
-- EXPRESS OR IMPLIED WARRANTIES, INCLUDING, BUT NOT LIMITED TO,
-- THE IMPLIED WARRANTIES OF MERCHANTABILITY AND FITNESS FOR A
-- PARTICULAR PURPOSE ARE DISCLAIMED. IN NO EVENT SHALL THE
-- ZPU PROJECT OR CONTRIBUTORS BE LIABLE FOR ANY DIRECT,
-- INDIRECT, INCIDENTAL, SPECIAL, EXEMPLARY, OR CONSEQUENTIAL DAMAGES
-- (INCLUDING, BUT NOT LIMITED TO, PROCUREMENT OF SUBSTITUTE GOODS
-- OR SERVICES; LOSS OF USE, DATA, OR PROFITS; OR BUSINESS INTERRUPTION)
-- HOWEVER CAUSED AND ON ANY THEORY OF LIABILITY, WHETHER IN CONTRACT,
-- STRICT LIABILITY, OR TORT (INCLUDING NEGLIGENCE OR OTHERWISE)
-- ARISING IN ANY WAY OUT OF THE USE OF THIS SOFTWARE, EVEN IF
-- ADVISED OF THE POSSIBILITY OF SUCH DAMAGE.
-- 
-- The views and conclusions contained in the software and documentation
-- are those of the authors and should not be interpreted as representing
-- official policies, either expressed or implied, of the ZPU Project.

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;


library work;
use work.zpu_config.all;
use work.zpupkg.all;

entity Dhrystone_min_ROM is
generic
	(
		maxAddrBitBRAM : integer := maxAddrBitBRAMLimit -- Specify your actual ROM size to save LEs and unnecessary block RAM usage.
	);
port (
	clk : in std_logic;
	areset : in std_logic := '0';
	from_zpu : in ZPU_ToROM;
	to_zpu : out ZPU_FromROM
);
end Dhrystone_min_ROM;

architecture arch of Dhrystone_min_ROM is

type ram_type is array(natural range 0 to ((2**(maxAddrBitBRAM+1))/4)-1) of std_logic_vector(wordSize-1 downto 0);

shared variable ram : ram_type :=
(
     0 => x"0b0b0b88",
     1 => x"dd040000",
     2 => x"00000000",
     3 => x"00000000",
     4 => x"00000000",
     5 => x"00000000",
     6 => x"00000000",
     7 => x"00000000",
     8 => x"88088c08",
     9 => x"90080b0b",
    10 => x"0b88e708",
    11 => x"2d900c8c",
    12 => x"0c880c04",
    13 => x"00000000",
    14 => x"00000000",
    15 => x"00000000",
    16 => x"71fd0608",
    17 => x"72830609",
    18 => x"81058205",
    19 => x"832b2a83",
    20 => x"ffff0652",
    21 => x"04000000",
    22 => x"00000000",
    23 => x"00000000",
    24 => x"71fd0608",
    25 => x"83ffff73",
    26 => x"83060981",
    27 => x"05820583",
    28 => x"2b2b0906",
    29 => x"7383ffff",
    30 => x"0b0b0b0b",
    31 => x"83a50400",
    32 => x"72098105",
    33 => x"72057373",
    34 => x"09060906",
    35 => x"73097306",
    36 => x"070a8106",
    37 => x"53510400",
    38 => x"00000000",
    39 => x"00000000",
    40 => x"72722473",
    41 => x"732e0753",
    42 => x"51040000",
    43 => x"00000000",
    44 => x"00000000",
    45 => x"00000000",
    46 => x"00000000",
    47 => x"00000000",
    48 => x"71737109",
    49 => x"71068106",
    50 => x"09810572",
    51 => x"0a100a72",
    52 => x"0a100a31",
    53 => x"050a8106",
    54 => x"51515351",
    55 => x"04000000",
    56 => x"72722673",
    57 => x"732e0753",
    58 => x"51040000",
    59 => x"00000000",
    60 => x"00000000",
    61 => x"00000000",
    62 => x"00000000",
    63 => x"00000000",
    64 => x"00000000",
    65 => x"00000000",
    66 => x"00000000",
    67 => x"00000000",
    68 => x"00000000",
    69 => x"00000000",
    70 => x"00000000",
    71 => x"00000000",
    72 => x"0b0b0b88",
    73 => x"ba040000",
    74 => x"00000000",
    75 => x"00000000",
    76 => x"00000000",
    77 => x"00000000",
    78 => x"00000000",
    79 => x"00000000",
    80 => x"720a722b",
    81 => x"0a535104",
    82 => x"00000000",
    83 => x"00000000",
    84 => x"00000000",
    85 => x"00000000",
    86 => x"00000000",
    87 => x"00000000",
    88 => x"72729f06",
    89 => x"0981050b",
    90 => x"0b0b889f",
    91 => x"05040000",
    92 => x"00000000",
    93 => x"00000000",
    94 => x"00000000",
    95 => x"00000000",
    96 => x"72722aff",
    97 => x"739f062a",
    98 => x"0974090a",
    99 => x"8106ff05",
   100 => x"06075351",
   101 => x"04000000",
   102 => x"00000000",
   103 => x"00000000",
   104 => x"71715351",
   105 => x"04067383",
   106 => x"06098105",
   107 => x"8205832b",
   108 => x"0b2b0772",
   109 => x"fc060c51",
   110 => x"51040000",
   111 => x"00000000",
   112 => x"72098105",
   113 => x"72050970",
   114 => x"81050906",
   115 => x"0a810653",
   116 => x"51040000",
   117 => x"00000000",
   118 => x"00000000",
   119 => x"00000000",
   120 => x"72098105",
   121 => x"72050970",
   122 => x"81050906",
   123 => x"0a098106",
   124 => x"53510400",
   125 => x"00000000",
   126 => x"00000000",
   127 => x"00000000",
   128 => x"71098105",
   129 => x"52040000",
   130 => x"00000000",
   131 => x"00000000",
   132 => x"00000000",
   133 => x"00000000",
   134 => x"00000000",
   135 => x"00000000",
   136 => x"72720981",
   137 => x"05055351",
   138 => x"04000000",
   139 => x"00000000",
   140 => x"00000000",
   141 => x"00000000",
   142 => x"00000000",
   143 => x"00000000",
   144 => x"72097206",
   145 => x"73730906",
   146 => x"07535104",
   147 => x"00000000",
   148 => x"00000000",
   149 => x"00000000",
   150 => x"00000000",
   151 => x"00000000",
   152 => x"71fc0608",
   153 => x"72830609",
   154 => x"81058305",
   155 => x"1010102a",
   156 => x"81ff0652",
   157 => x"04000000",
   158 => x"00000000",
   159 => x"00000000",
   160 => x"71fc0608",
   161 => x"0b0b0b9f",
   162 => x"a8738306",
   163 => x"10100508",
   164 => x"060b0b0b",
   165 => x"88a20400",
   166 => x"00000000",
   167 => x"00000000",
   168 => x"88088c08",
   169 => x"90087575",
   170 => x"0b0b0b98",
   171 => x"9c2d5050",
   172 => x"88085690",
   173 => x"0c8c0c88",
   174 => x"0c510400",
   175 => x"00000000",
   176 => x"88088c08",
   177 => x"90087575",
   178 => x"0b0b0b99",
   179 => x"ce2d5050",
   180 => x"88085690",
   181 => x"0c8c0c88",
   182 => x"0c510400",
   183 => x"00000000",
   184 => x"72097081",
   185 => x"0509060a",
   186 => x"8106ff05",
   187 => x"70547106",
   188 => x"73097274",
   189 => x"05ff0506",
   190 => x"07515151",
   191 => x"04000000",
   192 => x"72097081",
   193 => x"0509060a",
   194 => x"098106ff",
   195 => x"05705471",
   196 => x"06730972",
   197 => x"7405ff05",
   198 => x"06075151",
   199 => x"51040000",
   200 => x"05ff0504",
   201 => x"00000000",
   202 => x"00000000",
   203 => x"00000000",
   204 => x"00000000",
   205 => x"00000000",
   206 => x"00000000",
   207 => x"00000000",
   208 => x"04000000",
   209 => x"00000000",
   210 => x"00000000",
   211 => x"00000000",
   212 => x"00000000",
   213 => x"00000000",
   214 => x"00000000",
   215 => x"00000000",
   216 => x"71810552",
   217 => x"04000000",
   218 => x"00000000",
   219 => x"00000000",
   220 => x"00000000",
   221 => x"00000000",
   222 => x"00000000",
   223 => x"00000000",
   224 => x"00000000",
   225 => x"00000000",
   226 => x"00000000",
   227 => x"00000000",
   228 => x"00000000",
   229 => x"00000000",
   230 => x"00000000",
   231 => x"00000000",
   232 => x"02840572",
   233 => x"10100552",
   234 => x"04000000",
   235 => x"00000000",
   236 => x"00000000",
   237 => x"00000000",
   238 => x"00000000",
   239 => x"00000000",
   240 => x"00000000",
   241 => x"00000000",
   242 => x"00000000",
   243 => x"00000000",
   244 => x"00000000",
   245 => x"00000000",
   246 => x"00000000",
   247 => x"00000000",
   248 => x"717105ff",
   249 => x"05715351",
   250 => x"020d0400",
   251 => x"00000000",
   252 => x"00000000",
   253 => x"00000000",
   254 => x"00000000",
   255 => x"00000000",
   256 => x"10101010",
   257 => x"10101010",
   258 => x"10101010",
   259 => x"10101010",
   260 => x"10101010",
   261 => x"10101010",
   262 => x"10101010",
   263 => x"10101053",
   264 => x"51047381",
   265 => x"ff067383",
   266 => x"06098105",
   267 => x"83051010",
   268 => x"102b0772",
   269 => x"fc060c51",
   270 => x"51047272",
   271 => x"80728106",
   272 => x"ff050972",
   273 => x"06057110",
   274 => x"52720a10",
   275 => x"0a5372ed",
   276 => x"38515153",
   277 => x"51040000",
   278 => x"800488da",
   279 => x"0488da0b",
   280 => x"8efb0404",
   281 => x"00000000",
   282 => x"000463f0",
   283 => x"3d0d933d",
   284 => x"0b0b0ba4",
   285 => x"d05b5d80",
   286 => x"7d708405",
   287 => x"5f087140",
   288 => x"40587e70",
   289 => x"84054008",
   290 => x"57805976",
   291 => x"982a7788",
   292 => x"2b585574",
   293 => x"802e82af",
   294 => x"387d802e",
   295 => x"b738805e",
   296 => x"7480e42e",
   297 => x"81983874",
   298 => x"80e42680",
   299 => x"d8387480",
   300 => x"e32eb738",
   301 => x"a55182a0",
   302 => x"3f745182",
   303 => x"9b3f8218",
   304 => x"58811959",
   305 => x"837925c3",
   306 => x"3874ffb6",
   307 => x"387f880c",
   308 => x"923d0d04",
   309 => x"74a52e09",
   310 => x"81069738",
   311 => x"810b811a",
   312 => x"5a5e8379",
   313 => x"25ffa438",
   314 => x"e0397c84",
   315 => x"1e710857",
   316 => x"5e567451",
   317 => x"81e23f81",
   318 => x"18811a5a",
   319 => x"58837925",
   320 => x"ff8938c5",
   321 => x"397480f3",
   322 => x"2e098106",
   323 => x"ffa6387c",
   324 => x"841e7108",
   325 => x"70545c5e",
   326 => x"5481dc3f",
   327 => x"800bff11",
   328 => x"55538073",
   329 => x"25ff9a38",
   330 => x"79708105",
   331 => x"5b337052",
   332 => x"5581a53f",
   333 => x"811874ff",
   334 => x"16565458",
   335 => x"e5397c84",
   336 => x"1e71080b",
   337 => x"0b0ba4d0",
   338 => x"0b0b0b0b",
   339 => x"a4806240",
   340 => x"5a5f565e",
   341 => x"53807424",
   342 => x"80f43873",
   343 => x"b138b00b",
   344 => x"0b0b0ba4",
   345 => x"80348116",
   346 => x"56ff1656",
   347 => x"75337c70",
   348 => x"81055e34",
   349 => x"811b5b75",
   350 => x"0b0b0ba4",
   351 => x"802e0981",
   352 => x"06e73880",
   353 => x"7c347aff",
   354 => x"115553ff",
   355 => x"95398a74",
   356 => x"369fb805",
   357 => x"53723376",
   358 => x"70810558",
   359 => x"348a7435",
   360 => x"5473eb38",
   361 => x"750b0b0b",
   362 => x"a4802ed7",
   363 => x"38ff1656",
   364 => x"75337c70",
   365 => x"81055e34",
   366 => x"811b5b75",
   367 => x"0b0b0ba4",
   368 => x"802ec038",
   369 => x"ffa33977",
   370 => x"880c923d",
   371 => x"0d04ad51",
   372 => x"873f7330",
   373 => x"54ff8439",
   374 => x"ff3d0d73",
   375 => x"52c00870",
   376 => x"882a7081",
   377 => x"06515151",
   378 => x"70802ef1",
   379 => x"3871c00c",
   380 => x"71880c83",
   381 => x"3d0d04fb",
   382 => x"3d0d8078",
   383 => x"57557570",
   384 => x"84055708",
   385 => x"53805472",
   386 => x"982a7388",
   387 => x"2b545271",
   388 => x"802ea238",
   389 => x"c0087088",
   390 => x"2a708106",
   391 => x"51515170",
   392 => x"802ef138",
   393 => x"71c00c81",
   394 => x"15811555",
   395 => x"55837425",
   396 => x"d63871ca",
   397 => x"3874880c",
   398 => x"873d0d04",
   399 => x"c808880c",
   400 => x"04803d0d",
   401 => x"80c10b80",
   402 => x"f49c3480",
   403 => x"0b80f6b4",
   404 => x"0c70880c",
   405 => x"823d0d04",
   406 => x"ff3d0d80",
   407 => x"0b80f49c",
   408 => x"33525270",
   409 => x"80c12e99",
   410 => x"387180f6",
   411 => x"b4080780",
   412 => x"f6b40c80",
   413 => x"c20b80f4",
   414 => x"a0347088",
   415 => x"0c833d0d",
   416 => x"04810b80",
   417 => x"f6b40807",
   418 => x"80f6b40c",
   419 => x"80c20b80",
   420 => x"f4a03470",
   421 => x"880c833d",
   422 => x"0d04fd3d",
   423 => x"0d757008",
   424 => x"8a055353",
   425 => x"80f49c33",
   426 => x"517080c1",
   427 => x"2e8b3873",
   428 => x"f3387088",
   429 => x"0c853d0d",
   430 => x"04ff1270",
   431 => x"80f49808",
   432 => x"31740c88",
   433 => x"0c853d0d",
   434 => x"04fc3d0d",
   435 => x"80f4c408",
   436 => x"5574802e",
   437 => x"8c387675",
   438 => x"08710c80",
   439 => x"f4c40856",
   440 => x"548c1553",
   441 => x"80f49808",
   442 => x"528a5188",
   443 => x"9c3f7388",
   444 => x"0c863d0d",
   445 => x"04fb3d0d",
   446 => x"77700856",
   447 => x"56b05380",
   448 => x"f4c40852",
   449 => x"74518ef2",
   450 => x"3f850b8c",
   451 => x"170c850b",
   452 => x"8c160c75",
   453 => x"08750c80",
   454 => x"f4c40854",
   455 => x"73802e8a",
   456 => x"38730875",
   457 => x"0c80f4c4",
   458 => x"08548c14",
   459 => x"5380f498",
   460 => x"08528a51",
   461 => x"87d33f84",
   462 => x"1508ad38",
   463 => x"860b8c16",
   464 => x"0c881552",
   465 => x"88160851",
   466 => x"86df3f80",
   467 => x"f4c40870",
   468 => x"08760c54",
   469 => x"8c157054",
   470 => x"548a5273",
   471 => x"085187a9",
   472 => x"3f73880c",
   473 => x"873d0d04",
   474 => x"750854b0",
   475 => x"53735275",
   476 => x"518e873f",
   477 => x"73880c87",
   478 => x"3d0d04f3",
   479 => x"3d0d80f3",
   480 => x"b00b80f3",
   481 => x"e40c80f3",
   482 => x"e80b80f4",
   483 => x"c40c80f3",
   484 => x"b00b80f3",
   485 => x"e80c800b",
   486 => x"80f3e80b",
   487 => x"84050c82",
   488 => x"0b80f3e8",
   489 => x"0b88050c",
   490 => x"a80b80f3",
   491 => x"e80b8c05",
   492 => x"0c9f539f",
   493 => x"cc5280f3",
   494 => x"f8518dbe",
   495 => x"3f9f539f",
   496 => x"ec5280f6",
   497 => x"94518db2",
   498 => x"3f8a0bb1",
   499 => x"fc0ca2cc",
   500 => x"51f9983f",
   501 => x"a08c51f9",
   502 => x"923fa2cc",
   503 => x"51f98c3f",
   504 => x"a3fc0880",
   505 => x"2e83e638",
   506 => x"a0bc51f8",
   507 => x"fe3fa2cc",
   508 => x"51f8f83f",
   509 => x"a3f80852",
   510 => x"a0e851f8",
   511 => x"ee3fc808",
   512 => x"70a59c0c",
   513 => x"56815880",
   514 => x"0ba3f808",
   515 => x"2582c438",
   516 => x"8c3d5b80",
   517 => x"c10b80f4",
   518 => x"9c34810b",
   519 => x"80f6b40c",
   520 => x"80c20b80",
   521 => x"f4a03482",
   522 => x"5c835a9f",
   523 => x"53a19852",
   524 => x"80f4a451",
   525 => x"8cc43f81",
   526 => x"5d800b80",
   527 => x"f4a45380",
   528 => x"f6945255",
   529 => x"86e73f88",
   530 => x"08752e09",
   531 => x"81068338",
   532 => x"81557480",
   533 => x"f6b40c7b",
   534 => x"70575574",
   535 => x"8325a038",
   536 => x"74101015",
   537 => x"fd055e8f",
   538 => x"3dfc0553",
   539 => x"83527551",
   540 => x"85973f81",
   541 => x"1c705d70",
   542 => x"57558375",
   543 => x"24e2387d",
   544 => x"547453a5",
   545 => x"a05280f4",
   546 => x"cc51858d",
   547 => x"3f80f4c4",
   548 => x"08700857",
   549 => x"57b05376",
   550 => x"5275518b",
   551 => x"dd3f850b",
   552 => x"8c180c85",
   553 => x"0b8c170c",
   554 => x"7608760c",
   555 => x"80f4c408",
   556 => x"5574802e",
   557 => x"8a387408",
   558 => x"760c80f4",
   559 => x"c408558c",
   560 => x"155380f4",
   561 => x"9808528a",
   562 => x"5184be3f",
   563 => x"84160883",
   564 => x"9e38860b",
   565 => x"8c170c88",
   566 => x"16528817",
   567 => x"085183c9",
   568 => x"3f80f4c4",
   569 => x"08700877",
   570 => x"0c578c16",
   571 => x"7054558a",
   572 => x"52740851",
   573 => x"84933f80",
   574 => x"c10b80f4",
   575 => x"a0335656",
   576 => x"757526a2",
   577 => x"3880c352",
   578 => x"755184f7",
   579 => x"3f88087d",
   580 => x"2e82af38",
   581 => x"81167081",
   582 => x"ff0680f4",
   583 => x"a0335257",
   584 => x"55747627",
   585 => x"e0387d7a",
   586 => x"7d293570",
   587 => x"5d8a0580",
   588 => x"f49c3380",
   589 => x"f4980859",
   590 => x"57557580",
   591 => x"c12e82c7",
   592 => x"3878f738",
   593 => x"811858a3",
   594 => x"f8087825",
   595 => x"fdc538a5",
   596 => x"9c0856c8",
   597 => x"087080f3",
   598 => x"e00c7077",
   599 => x"3170a598",
   600 => x"0c53a1b8",
   601 => x"525bf683",
   602 => x"3fa59808",
   603 => x"5680f776",
   604 => x"2580e038",
   605 => x"a3f80870",
   606 => x"7787e829",
   607 => x"35a5900c",
   608 => x"767187e8",
   609 => x"2935a594",
   610 => x"0c767184",
   611 => x"b9293580",
   612 => x"f4c80c5a",
   613 => x"a1c851f5",
   614 => x"d23fa590",
   615 => x"0852a1f8",
   616 => x"51f5c83f",
   617 => x"a28051f5",
   618 => x"c23fa594",
   619 => x"0852a1f8",
   620 => x"51f5b83f",
   621 => x"80f4c808",
   622 => x"52a2b051",
   623 => x"f5ad3fa2",
   624 => x"cc51f5a7",
   625 => x"3f800b88",
   626 => x"0c8f3d0d",
   627 => x"04a2d051",
   628 => x"fc9939a3",
   629 => x"8051f593",
   630 => x"3fa3b851",
   631 => x"f58d3fa2",
   632 => x"cc51f587",
   633 => x"3fa59808",
   634 => x"a3f80870",
   635 => x"7287e829",
   636 => x"35a5900c",
   637 => x"717187e8",
   638 => x"2935a594",
   639 => x"0c717184",
   640 => x"b9293580",
   641 => x"f4c80c5b",
   642 => x"56a1c851",
   643 => x"f4dd3fa5",
   644 => x"900852a1",
   645 => x"f851f4d3",
   646 => x"3fa28051",
   647 => x"f4cd3fa5",
   648 => x"940852a1",
   649 => x"f851f4c3",
   650 => x"3f80f4c8",
   651 => x"0852a2b0",
   652 => x"51f4b83f",
   653 => x"a2cc51f4",
   654 => x"b23f800b",
   655 => x"880c8f3d",
   656 => x"0d048f3d",
   657 => x"f8055280",
   658 => x"5180de3f",
   659 => x"9f53a3d8",
   660 => x"5280f4a4",
   661 => x"5188a33f",
   662 => x"777880f4",
   663 => x"980c8117",
   664 => x"7081ff06",
   665 => x"80f4a033",
   666 => x"5258565a",
   667 => x"fdb33976",
   668 => x"0856b053",
   669 => x"75527651",
   670 => x"88803f80",
   671 => x"c10b80f4",
   672 => x"a0335656",
   673 => x"fcfa39ff",
   674 => x"15707831",
   675 => x"7c0c5980",
   676 => x"59fdb139",
   677 => x"ff3d0d73",
   678 => x"82327030",
   679 => x"70720780",
   680 => x"25880c52",
   681 => x"52833d0d",
   682 => x"04fe3d0d",
   683 => x"74767153",
   684 => x"54527182",
   685 => x"2e833883",
   686 => x"5171812e",
   687 => x"9a388172",
   688 => x"269f3871",
   689 => x"822eb838",
   690 => x"71842ea9",
   691 => x"3870730c",
   692 => x"70880c84",
   693 => x"3d0d0480",
   694 => x"e40b80f4",
   695 => x"9808258b",
   696 => x"3880730c",
   697 => x"70880c84",
   698 => x"3d0d0483",
   699 => x"730c7088",
   700 => x"0c843d0d",
   701 => x"0482730c",
   702 => x"70880c84",
   703 => x"3d0d0481",
   704 => x"730c7088",
   705 => x"0c843d0d",
   706 => x"04803d0d",
   707 => x"74741482",
   708 => x"05710c88",
   709 => x"0c823d0d",
   710 => x"04f73d0d",
   711 => x"7b7d7f61",
   712 => x"85127082",
   713 => x"2b751170",
   714 => x"74717084",
   715 => x"05530c5a",
   716 => x"5a5d5b76",
   717 => x"0c7980f8",
   718 => x"180c7986",
   719 => x"12525758",
   720 => x"5a5a7676",
   721 => x"24993876",
   722 => x"b329822b",
   723 => x"79115153",
   724 => x"76737084",
   725 => x"05550c81",
   726 => x"14547574",
   727 => x"25f23876",
   728 => x"81cc2919",
   729 => x"fc110881",
   730 => x"05fc120c",
   731 => x"7a197008",
   732 => x"9fa0130c",
   733 => x"5856850b",
   734 => x"80f4980c",
   735 => x"75880c8b",
   736 => x"3d0d04fe",
   737 => x"3d0d0293",
   738 => x"05335180",
   739 => x"02840597",
   740 => x"05335452",
   741 => x"70732e88",
   742 => x"3871880c",
   743 => x"843d0d04",
   744 => x"7080f49c",
   745 => x"34810b88",
   746 => x"0c843d0d",
   747 => x"04f83d0d",
   748 => x"7a7c5956",
   749 => x"820b8319",
   750 => x"55557416",
   751 => x"70337533",
   752 => x"5b515372",
   753 => x"792e80c6",
   754 => x"3880c10b",
   755 => x"81168116",
   756 => x"56565782",
   757 => x"7525e338",
   758 => x"ffa91770",
   759 => x"81ff0655",
   760 => x"59738226",
   761 => x"83388755",
   762 => x"81537680",
   763 => x"d22e9838",
   764 => x"77527551",
   765 => x"869d3f80",
   766 => x"53728808",
   767 => x"25893887",
   768 => x"1580f498",
   769 => x"0c815372",
   770 => x"880c8a3d",
   771 => x"0d047280",
   772 => x"f49c3482",
   773 => x"7525ffa2",
   774 => x"38ffbd39",
   775 => x"94080294",
   776 => x"0cf93d0d",
   777 => x"800b9408",
   778 => x"fc050c94",
   779 => x"08880508",
   780 => x"8025ab38",
   781 => x"94088805",
   782 => x"08309408",
   783 => x"88050c80",
   784 => x"0b9408f4",
   785 => x"050c9408",
   786 => x"fc050888",
   787 => x"38810b94",
   788 => x"08f4050c",
   789 => x"9408f405",
   790 => x"089408fc",
   791 => x"050c9408",
   792 => x"8c050880",
   793 => x"25ab3894",
   794 => x"088c0508",
   795 => x"3094088c",
   796 => x"050c800b",
   797 => x"9408f005",
   798 => x"0c9408fc",
   799 => x"05088838",
   800 => x"810b9408",
   801 => x"f0050c94",
   802 => x"08f00508",
   803 => x"9408fc05",
   804 => x"0c805394",
   805 => x"088c0508",
   806 => x"52940888",
   807 => x"05085181",
   808 => x"a73f8808",
   809 => x"709408f8",
   810 => x"050c5494",
   811 => x"08fc0508",
   812 => x"802e8c38",
   813 => x"9408f805",
   814 => x"08309408",
   815 => x"f8050c94",
   816 => x"08f80508",
   817 => x"70880c54",
   818 => x"893d0d94",
   819 => x"0c049408",
   820 => x"02940cfb",
   821 => x"3d0d800b",
   822 => x"9408fc05",
   823 => x"0c940888",
   824 => x"05088025",
   825 => x"93389408",
   826 => x"88050830",
   827 => x"94088805",
   828 => x"0c810b94",
   829 => x"08fc050c",
   830 => x"94088c05",
   831 => x"0880258c",
   832 => x"3894088c",
   833 => x"05083094",
   834 => x"088c050c",
   835 => x"81539408",
   836 => x"8c050852",
   837 => x"94088805",
   838 => x"0851ad3f",
   839 => x"88087094",
   840 => x"08f8050c",
   841 => x"549408fc",
   842 => x"0508802e",
   843 => x"8c389408",
   844 => x"f8050830",
   845 => x"9408f805",
   846 => x"0c9408f8",
   847 => x"05087088",
   848 => x"0c54873d",
   849 => x"0d940c04",
   850 => x"94080294",
   851 => x"0cfd3d0d",
   852 => x"810b9408",
   853 => x"fc050c80",
   854 => x"0b9408f8",
   855 => x"050c9408",
   856 => x"8c050894",
   857 => x"08880508",
   858 => x"27ac3894",
   859 => x"08fc0508",
   860 => x"802ea338",
   861 => x"800b9408",
   862 => x"8c050824",
   863 => x"99389408",
   864 => x"8c050810",
   865 => x"94088c05",
   866 => x"0c9408fc",
   867 => x"05081094",
   868 => x"08fc050c",
   869 => x"c9399408",
   870 => x"fc050880",
   871 => x"2e80c938",
   872 => x"94088c05",
   873 => x"08940888",
   874 => x"050826a1",
   875 => x"38940888",
   876 => x"05089408",
   877 => x"8c050831",
   878 => x"94088805",
   879 => x"0c9408f8",
   880 => x"05089408",
   881 => x"fc050807",
   882 => x"9408f805",
   883 => x"0c9408fc",
   884 => x"0508812a",
   885 => x"9408fc05",
   886 => x"0c94088c",
   887 => x"0508812a",
   888 => x"94088c05",
   889 => x"0cffaf39",
   890 => x"94089005",
   891 => x"08802e8f",
   892 => x"38940888",
   893 => x"05087094",
   894 => x"08f4050c",
   895 => x"518d3994",
   896 => x"08f80508",
   897 => x"709408f4",
   898 => x"050c5194",
   899 => x"08f40508",
   900 => x"880c853d",
   901 => x"0d940c04",
   902 => x"94080294",
   903 => x"0cff3d0d",
   904 => x"800b9408",
   905 => x"fc050c94",
   906 => x"08880508",
   907 => x"8106ff11",
   908 => x"70097094",
   909 => x"088c0508",
   910 => x"069408fc",
   911 => x"05081194",
   912 => x"08fc050c",
   913 => x"94088805",
   914 => x"08812a94",
   915 => x"0888050c",
   916 => x"94088c05",
   917 => x"08109408",
   918 => x"8c050c51",
   919 => x"51515194",
   920 => x"08880508",
   921 => x"802e8438",
   922 => x"ffbd3994",
   923 => x"08fc0508",
   924 => x"70880c51",
   925 => x"833d0d94",
   926 => x"0c04fc3d",
   927 => x"0d767079",
   928 => x"7b555555",
   929 => x"558f7227",
   930 => x"8c387275",
   931 => x"07830651",
   932 => x"70802ea7",
   933 => x"38ff1252",
   934 => x"71ff2e98",
   935 => x"38727081",
   936 => x"05543374",
   937 => x"70810556",
   938 => x"34ff1252",
   939 => x"71ff2e09",
   940 => x"8106ea38",
   941 => x"74880c86",
   942 => x"3d0d0474",
   943 => x"51727084",
   944 => x"05540871",
   945 => x"70840553",
   946 => x"0c727084",
   947 => x"05540871",
   948 => x"70840553",
   949 => x"0c727084",
   950 => x"05540871",
   951 => x"70840553",
   952 => x"0c727084",
   953 => x"05540871",
   954 => x"70840553",
   955 => x"0cf01252",
   956 => x"718f26c9",
   957 => x"38837227",
   958 => x"95387270",
   959 => x"84055408",
   960 => x"71708405",
   961 => x"530cfc12",
   962 => x"52718326",
   963 => x"ed387054",
   964 => x"ff8339fb",
   965 => x"3d0d7779",
   966 => x"70720783",
   967 => x"06535452",
   968 => x"70933871",
   969 => x"73730854",
   970 => x"56547173",
   971 => x"082e80c4",
   972 => x"38737554",
   973 => x"52713370",
   974 => x"81ff0652",
   975 => x"5470802e",
   976 => x"9d387233",
   977 => x"5570752e",
   978 => x"09810695",
   979 => x"38811281",
   980 => x"14713370",
   981 => x"81ff0654",
   982 => x"56545270",
   983 => x"e5387233",
   984 => x"557381ff",
   985 => x"067581ff",
   986 => x"06717131",
   987 => x"880c5252",
   988 => x"873d0d04",
   989 => x"710970f7",
   990 => x"fbfdff14",
   991 => x"0670f884",
   992 => x"82818006",
   993 => x"51515170",
   994 => x"97388414",
   995 => x"84167108",
   996 => x"54565471",
   997 => x"75082edc",
   998 => x"38737554",
   999 => x"52ff9639",
  1000 => x"800b880c",
  1001 => x"873d0d04",
  1002 => x"00ffffff",
  1003 => x"ff00ffff",
  1004 => x"ffff00ff",
  1005 => x"ffffff00",
  1006 => x"30313233",
  1007 => x"34353637",
  1008 => x"38394142",
  1009 => x"43444546",
  1010 => x"00000000",
  1011 => x"44485259",
  1012 => x"53544f4e",
  1013 => x"45205052",
  1014 => x"4f475241",
  1015 => x"4d2c2053",
  1016 => x"4f4d4520",
  1017 => x"53545249",
  1018 => x"4e470000",
  1019 => x"44485259",
  1020 => x"53544f4e",
  1021 => x"45205052",
  1022 => x"4f475241",
  1023 => x"4d2c2031",
  1024 => x"27535420",
  1025 => x"53545249",
  1026 => x"4e470000",
  1027 => x"44687279",
  1028 => x"73746f6e",
  1029 => x"65204265",
  1030 => x"6e63686d",
  1031 => x"61726b2c",
  1032 => x"20566572",
  1033 => x"73696f6e",
  1034 => x"20322e31",
  1035 => x"20284c61",
  1036 => x"6e677561",
  1037 => x"67653a20",
  1038 => x"43290a00",
  1039 => x"50726f67",
  1040 => x"72616d20",
  1041 => x"636f6d70",
  1042 => x"696c6564",
  1043 => x"20776974",
  1044 => x"68202772",
  1045 => x"65676973",
  1046 => x"74657227",
  1047 => x"20617474",
  1048 => x"72696275",
  1049 => x"74650a00",
  1050 => x"45786563",
  1051 => x"7574696f",
  1052 => x"6e207374",
  1053 => x"61727473",
  1054 => x"2c202564",
  1055 => x"2072756e",
  1056 => x"73207468",
  1057 => x"726f7567",
  1058 => x"68204468",
  1059 => x"72797374",
  1060 => x"6f6e650a",
  1061 => x"00000000",
  1062 => x"44485259",
  1063 => x"53544f4e",
  1064 => x"45205052",
  1065 => x"4f475241",
  1066 => x"4d2c2032",
  1067 => x"274e4420",
  1068 => x"53545249",
  1069 => x"4e470000",
  1070 => x"55736572",
  1071 => x"2074696d",
  1072 => x"653a2025",
  1073 => x"640a0000",
  1074 => x"4d696372",
  1075 => x"6f736563",
  1076 => x"6f6e6473",
  1077 => x"20666f72",
  1078 => x"206f6e65",
  1079 => x"2072756e",
  1080 => x"20746872",
  1081 => x"6f756768",
  1082 => x"20446872",
  1083 => x"7973746f",
  1084 => x"6e653a20",
  1085 => x"00000000",
  1086 => x"2564200a",
  1087 => x"00000000",
  1088 => x"44687279",
  1089 => x"73746f6e",
  1090 => x"65732070",
  1091 => x"65722053",
  1092 => x"65636f6e",
  1093 => x"643a2020",
  1094 => x"20202020",
  1095 => x"20202020",
  1096 => x"20202020",
  1097 => x"20202020",
  1098 => x"20202020",
  1099 => x"00000000",
  1100 => x"56415820",
  1101 => x"4d495053",
  1102 => x"20726174",
  1103 => x"696e6720",
  1104 => x"2a203130",
  1105 => x"3030203d",
  1106 => x"20256420",
  1107 => x"0a000000",
  1108 => x"50726f67",
  1109 => x"72616d20",
  1110 => x"636f6d70",
  1111 => x"696c6564",
  1112 => x"20776974",
  1113 => x"686f7574",
  1114 => x"20277265",
  1115 => x"67697374",
  1116 => x"65722720",
  1117 => x"61747472",
  1118 => x"69627574",
  1119 => x"650a0000",
  1120 => x"4d656173",
  1121 => x"75726564",
  1122 => x"2074696d",
  1123 => x"6520746f",
  1124 => x"6f20736d",
  1125 => x"616c6c20",
  1126 => x"746f206f",
  1127 => x"62746169",
  1128 => x"6e206d65",
  1129 => x"616e696e",
  1130 => x"6766756c",
  1131 => x"20726573",
  1132 => x"756c7473",
  1133 => x"0a000000",
  1134 => x"506c6561",
  1135 => x"73652069",
  1136 => x"6e637265",
  1137 => x"61736520",
  1138 => x"6e756d62",
  1139 => x"6572206f",
  1140 => x"66207275",
  1141 => x"6e730a00",
  1142 => x"44485259",
  1143 => x"53544f4e",
  1144 => x"45205052",
  1145 => x"4f475241",
  1146 => x"4d2c2033",
  1147 => x"27524420",
  1148 => x"53545249",
  1149 => x"4e470000",
  1150 => x"000061a8",
  1151 => x"00000000",
	others => x"00000000"
);

begin

process (clk)
begin
	if (clk'event and clk = '1') then
		if (from_zpu.memAWriteEnable = '1') and (from_zpu.memBWriteEnable = '1') and (from_zpu.memAAddr=from_zpu.memBAddr) and (from_zpu.memAWrite/=from_zpu.memBWrite) then
			report "write collision" severity failure;
		end if;
	
		if (from_zpu.memAWriteEnable = '1') then
			ram(to_integer(unsigned(from_zpu.memAAddr(maxAddrBitBRAM downto 2)))) := from_zpu.memAWrite;
			to_zpu.memARead <= from_zpu.memAWrite;
		else
			to_zpu.memARead <= ram(to_integer(unsigned(from_zpu.memAAddr(maxAddrBitBRAM downto 2))));
		end if;
	end if;
end process;

process (clk)
begin
	if (clk'event and clk = '1') then
		if (from_zpu.memBWriteEnable = '1') then
			ram(to_integer(unsigned(from_zpu.memBAddr(maxAddrBitBRAM downto 2)))) := from_zpu.memBWrite;
			to_zpu.memBRead <= from_zpu.memBWrite;
		else
			to_zpu.memBRead <= ram(to_integer(unsigned(from_zpu.memBAddr(maxAddrBitBRAM downto 2))));
		end if;
	end if;
end process;


end arch;

