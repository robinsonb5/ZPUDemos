-- ZPU
--
-- Copyright 2004-2008 oharboe - �yvind Harboe - oyvind.harboe@zylin.com
-- Modified by Alastair M. Robinson for the ZPUFlex project.
--
-- The FreeBSD license
-- 
-- Redistribution and use in source and binary forms, with or without
-- modification, are permitted provided that the following conditions
-- are met:
-- 
-- 1. Redistributions of source code must retain the above copyright
--    notice, this list of conditions and the following disclaimer.
-- 2. Redistributions in binary form must reproduce the above
--    copyright notice, this list of conditions and the following
--    disclaimer in the documentation and/or other materials
--    provided with the distribution.
-- 
-- THIS SOFTWARE IS PROVIDED BY THE ZPU PROJECT ``AS IS'' AND ANY
-- EXPRESS OR IMPLIED WARRANTIES, INCLUDING, BUT NOT LIMITED TO,
-- THE IMPLIED WARRANTIES OF MERCHANTABILITY AND FITNESS FOR A
-- PARTICULAR PURPOSE ARE DISCLAIMED. IN NO EVENT SHALL THE
-- ZPU PROJECT OR CONTRIBUTORS BE LIABLE FOR ANY DIRECT,
-- INDIRECT, INCIDENTAL, SPECIAL, EXEMPLARY, OR CONSEQUENTIAL DAMAGES
-- (INCLUDING, BUT NOT LIMITED TO, PROCUREMENT OF SUBSTITUTE GOODS
-- OR SERVICES; LOSS OF USE, DATA, OR PROFITS; OR BUSINESS INTERRUPTION)
-- HOWEVER CAUSED AND ON ANY THEORY OF LIABILITY, WHETHER IN CONTRACT,
-- STRICT LIABILITY, OR TORT (INCLUDING NEGLIGENCE OR OTHERWISE)
-- ARISING IN ANY WAY OUT OF THE USE OF THIS SOFTWARE, EVEN IF
-- ADVISED OF THE POSSIBILITY OF SUCH DAMAGE.
-- 
-- The views and conclusions contained in the software and documentation
-- are those of the authors and should not be interpreted as representing
-- official policies, either expressed or implied, of the ZPU Project.

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;


library work;
use work.zpu_config.all;
use work.zpupkg.all;

entity SDBootstrap_ROM is
generic
	(
		maxAddrBitBRAM : integer := maxAddrBitBRAMLimit -- Specify your actual ROM size to save LEs and unnecessary block RAM usage.
	);
port (
	clk : in std_logic;
	areset : in std_logic := '0';
	from_zpu : in ZPU_ToROM;
	to_zpu : out ZPU_FromROM
);
end SDBootstrap_ROM;

architecture arch of SDBootstrap_ROM is

type ram_type is array(natural range 0 to ((2**(maxAddrBitBRAM+1))/4)-1) of std_logic_vector(wordSize-1 downto 0);

shared variable ram : ram_type :=
(
     0 => x"84808080",
     1 => x"ee040000",
     2 => x"00000000",
     3 => x"84808080",
     4 => x"88080d80",
     5 => x"04848080",
     6 => x"80950471",
     7 => x"fd060872",
     8 => x"83060981",
     9 => x"05820583",
    10 => x"2b2a83ff",
    11 => x"ff065204",
    12 => x"71fc0608",
    13 => x"72830609",
    14 => x"81058305",
    15 => x"1010102a",
    16 => x"81ff0652",
    17 => x"0471fc06",
    18 => x"08848080",
    19 => x"a1ec7383",
    20 => x"06101005",
    21 => x"08067381",
    22 => x"ff067383",
    23 => x"06098105",
    24 => x"83051010",
    25 => x"102b0772",
    26 => x"fc060c51",
    27 => x"51040284",
    28 => x"05848080",
    29 => x"80880c84",
    30 => x"80808095",
    31 => x"0b848080",
    32 => x"8ec50400",
    33 => x"02ec050d",
    34 => x"76538055",
    35 => x"7275258e",
    36 => x"38ad5184",
    37 => x"808084b2",
    38 => x"2d720981",
    39 => x"05537280",
    40 => x"2ebe3887",
    41 => x"54729c2a",
    42 => x"73842b54",
    43 => x"5271802e",
    44 => x"83388155",
    45 => x"8972258a",
    46 => x"38b71252",
    47 => x"84808081",
    48 => x"c504b012",
    49 => x"5274802e",
    50 => x"89387151",
    51 => x"84808084",
    52 => x"b22dff14",
    53 => x"54738025",
    54 => x"cc388480",
    55 => x"8081e804",
    56 => x"b0518480",
    57 => x"8084b22d",
    58 => x"800b83ff",
    59 => x"e0800c02",
    60 => x"94050d04",
    61 => x"02c0050d",
    62 => x"0280c405",
    63 => x"57807078",
    64 => x"7084055a",
    65 => x"0872415f",
    66 => x"5d587c70",
    67 => x"84055e08",
    68 => x"5a805b79",
    69 => x"982a7a88",
    70 => x"2b5b5675",
    71 => x"8938775f",
    72 => x"84808084",
    73 => x"a6047d80",
    74 => x"2e81d338",
    75 => x"805e7580",
    76 => x"e42e8a38",
    77 => x"7580f82e",
    78 => x"09810689",
    79 => x"38768418",
    80 => x"71085e58",
    81 => x"547580e4",
    82 => x"2ea63875",
    83 => x"80e4268e",
    84 => x"387580e3",
    85 => x"2e80d938",
    86 => x"84808083",
    87 => x"be047580",
    88 => x"f32eb538",
    89 => x"7580f82e",
    90 => x"8f388480",
    91 => x"8083be04",
    92 => x"8a538480",
    93 => x"8082fa04",
    94 => x"905383ff",
    95 => x"e0e0527b",
    96 => x"51848080",
    97 => x"81842d83",
    98 => x"ffe08008",
    99 => x"83ffe0e0",
   100 => x"5a558480",
   101 => x"8083d704",
   102 => x"76841871",
   103 => x"0870545b",
   104 => x"58548480",
   105 => x"8084d62d",
   106 => x"80558480",
   107 => x"8083d704",
   108 => x"76841871",
   109 => x"08585854",
   110 => x"84808084",
   111 => x"8e04a551",
   112 => x"84808084",
   113 => x"b22d7551",
   114 => x"84808084",
   115 => x"b22d8218",
   116 => x"58848080",
   117 => x"84990474",
   118 => x"ff165654",
   119 => x"807425b9",
   120 => x"38787081",
   121 => x"055a8480",
   122 => x"8080b02d",
   123 => x"70525684",
   124 => x"808084b2",
   125 => x"2d811858",
   126 => x"84808083",
   127 => x"d70475a5",
   128 => x"2e098106",
   129 => x"8938815e",
   130 => x"84808084",
   131 => x"99047551",
   132 => x"84808084",
   133 => x"b22d8118",
   134 => x"58811b5b",
   135 => x"837b25fd",
   136 => x"f23875fd",
   137 => x"e5387e83",
   138 => x"ffe0800c",
   139 => x"0280c005",
   140 => x"0d0402f8",
   141 => x"050d7352",
   142 => x"c0087088",
   143 => x"2a708106",
   144 => x"51515170",
   145 => x"802ef138",
   146 => x"71c00c71",
   147 => x"83ffe080",
   148 => x"0c028805",
   149 => x"0d0402e8",
   150 => x"050d8078",
   151 => x"57557570",
   152 => x"84055708",
   153 => x"53805472",
   154 => x"982a7388",
   155 => x"2b545271",
   156 => x"802ea238",
   157 => x"c0087088",
   158 => x"2a708106",
   159 => x"51515170",
   160 => x"802ef138",
   161 => x"71c00c81",
   162 => x"15811555",
   163 => x"55837425",
   164 => x"d63871ca",
   165 => x"387483ff",
   166 => x"e0800c02",
   167 => x"98050d04",
   168 => x"02f4050d",
   169 => x"d45281ff",
   170 => x"720c7108",
   171 => x"5381ff72",
   172 => x"0c72882b",
   173 => x"83fe8006",
   174 => x"72087081",
   175 => x"ff065152",
   176 => x"5381ff72",
   177 => x"0c727107",
   178 => x"882b7208",
   179 => x"7081ff06",
   180 => x"51525381",
   181 => x"ff720c72",
   182 => x"7107882b",
   183 => x"72087081",
   184 => x"ff067207",
   185 => x"83ffe080",
   186 => x"0c525302",
   187 => x"8c050d04",
   188 => x"02f4050d",
   189 => x"74767181",
   190 => x"ff06d40c",
   191 => x"535383ff",
   192 => x"f1a00885",
   193 => x"3871892b",
   194 => x"5271982a",
   195 => x"d40c7190",
   196 => x"2a7081ff",
   197 => x"06d40c51",
   198 => x"71882a70",
   199 => x"81ff06d4",
   200 => x"0c517181",
   201 => x"ff06d40c",
   202 => x"72902a70",
   203 => x"81ff06d4",
   204 => x"0c51d408",
   205 => x"7081ff06",
   206 => x"515182b8",
   207 => x"bf527081",
   208 => x"ff2e0981",
   209 => x"06943881",
   210 => x"ff0bd40c",
   211 => x"d4087081",
   212 => x"ff06ff14",
   213 => x"54515171",
   214 => x"e5387083",
   215 => x"ffe0800c",
   216 => x"028c050d",
   217 => x"0402fc05",
   218 => x"0d81c751",
   219 => x"81ff0bd4",
   220 => x"0cff1151",
   221 => x"708025f4",
   222 => x"38028405",
   223 => x"0d0402f0",
   224 => x"050d8480",
   225 => x"8086e52d",
   226 => x"819c9f53",
   227 => x"805287fc",
   228 => x"80f75184",
   229 => x"808085f0",
   230 => x"2d83ffe0",
   231 => x"80085483",
   232 => x"ffe08008",
   233 => x"812e0981",
   234 => x"06ae3881",
   235 => x"ff0bd40c",
   236 => x"820a5284",
   237 => x"9c80e951",
   238 => x"84808085",
   239 => x"f02d83ff",
   240 => x"e080088e",
   241 => x"3881ff0b",
   242 => x"d40c7353",
   243 => x"84808087",
   244 => x"df048480",
   245 => x"8086e52d",
   246 => x"ff135372",
   247 => x"ffae3872",
   248 => x"83ffe080",
   249 => x"0c029005",
   250 => x"0d0402f4",
   251 => x"050d81ff",
   252 => x"0bd40c84",
   253 => x"8080a1fc",
   254 => x"51848080",
   255 => x"84d62d93",
   256 => x"53805287",
   257 => x"fc80c151",
   258 => x"84808085",
   259 => x"f02d83ff",
   260 => x"e080088e",
   261 => x"3881ff0b",
   262 => x"d40c8153",
   263 => x"84808088",
   264 => x"ae048480",
   265 => x"8086e52d",
   266 => x"ff135372",
   267 => x"d4387283",
   268 => x"ffe0800c",
   269 => x"028c050d",
   270 => x"0402f005",
   271 => x"0d848080",
   272 => x"86e52d83",
   273 => x"aa52849c",
   274 => x"80c85184",
   275 => x"808085f0",
   276 => x"2d83ffe0",
   277 => x"800883ff",
   278 => x"e0800853",
   279 => x"848080a2",
   280 => x"88525384",
   281 => x"808081f4",
   282 => x"2d72812e",
   283 => x"098106a9",
   284 => x"38848080",
   285 => x"85a02d83",
   286 => x"ffe08008",
   287 => x"83ffff06",
   288 => x"537283aa",
   289 => x"2ebb3883",
   290 => x"ffe08008",
   291 => x"52848080",
   292 => x"a2a05184",
   293 => x"808081f4",
   294 => x"2d848080",
   295 => x"87ea2d84",
   296 => x"808089b9",
   297 => x"04815484",
   298 => x"80808ae4",
   299 => x"04848080",
   300 => x"a2b85184",
   301 => x"808081f4",
   302 => x"2d805484",
   303 => x"80808ae4",
   304 => x"0481ff0b",
   305 => x"d40cb153",
   306 => x"84808086",
   307 => x"fe2d83ff",
   308 => x"e0800880",
   309 => x"2e80fe38",
   310 => x"805287fc",
   311 => x"80fa5184",
   312 => x"808085f0",
   313 => x"2d83ffe0",
   314 => x"800880d7",
   315 => x"3883ffe0",
   316 => x"80085284",
   317 => x"8080a2d4",
   318 => x"51848080",
   319 => x"81f42d81",
   320 => x"ff0bd40c",
   321 => x"d4087081",
   322 => x"ff067054",
   323 => x"848080a2",
   324 => x"e0535153",
   325 => x"84808081",
   326 => x"f42d81ff",
   327 => x"0bd40c81",
   328 => x"ff0bd40c",
   329 => x"81ff0bd4",
   330 => x"0c81ff0b",
   331 => x"d40c7286",
   332 => x"2a708106",
   333 => x"70565153",
   334 => x"72802ea8",
   335 => x"38848080",
   336 => x"89a50483",
   337 => x"ffe08008",
   338 => x"52848080",
   339 => x"a2d45184",
   340 => x"808081f4",
   341 => x"2d72822e",
   342 => x"fed338ff",
   343 => x"135372fe",
   344 => x"e7387254",
   345 => x"7383ffe0",
   346 => x"800c0290",
   347 => x"050d0402",
   348 => x"f4050d81",
   349 => x"0b83fff1",
   350 => x"a00cd008",
   351 => x"708f2a70",
   352 => x"81065151",
   353 => x"5372f338",
   354 => x"72d00c84",
   355 => x"808086e5",
   356 => x"2dd00870",
   357 => x"8f2a7081",
   358 => x"06515153",
   359 => x"72f33881",
   360 => x"0bd00c87",
   361 => x"53805284",
   362 => x"d480c051",
   363 => x"84808085",
   364 => x"f02d83ff",
   365 => x"e0800881",
   366 => x"2e973872",
   367 => x"822e0981",
   368 => x"06893880",
   369 => x"53848080",
   370 => x"8c8b04ff",
   371 => x"135372d5",
   372 => x"38848080",
   373 => x"88b92d83",
   374 => x"ffe08008",
   375 => x"83fff1a0",
   376 => x"0c815287",
   377 => x"fc80d051",
   378 => x"84808085",
   379 => x"f02d81ff",
   380 => x"0bd40cd0",
   381 => x"08708f2a",
   382 => x"70810651",
   383 => x"515372f3",
   384 => x"3872d00c",
   385 => x"81ff0bd4",
   386 => x"0c815372",
   387 => x"83ffe080",
   388 => x"0c028c05",
   389 => x"0d04800b",
   390 => x"83ffe080",
   391 => x"0c0402e0",
   392 => x"050d797b",
   393 => x"57578058",
   394 => x"81ff0bd4",
   395 => x"0cd00870",
   396 => x"8f2a7081",
   397 => x"06515154",
   398 => x"73f33882",
   399 => x"810bd00c",
   400 => x"81ff0bd4",
   401 => x"0c765287",
   402 => x"fc80d151",
   403 => x"84808085",
   404 => x"f02d80db",
   405 => x"c6df5583",
   406 => x"ffe08008",
   407 => x"802e9b38",
   408 => x"83ffe080",
   409 => x"08537652",
   410 => x"848080a2",
   411 => x"f0518480",
   412 => x"8081f42d",
   413 => x"8480808d",
   414 => x"d00481ff",
   415 => x"0bd40cd4",
   416 => x"087081ff",
   417 => x"06515473",
   418 => x"81fe2e09",
   419 => x"8106a538",
   420 => x"80ff5484",
   421 => x"808085a0",
   422 => x"2d83ffe0",
   423 => x"80087670",
   424 => x"8405580c",
   425 => x"ff145473",
   426 => x"8025e838",
   427 => x"81588480",
   428 => x"808dba04",
   429 => x"ff155574",
   430 => x"c13881ff",
   431 => x"0bd40cd0",
   432 => x"08708f2a",
   433 => x"70810651",
   434 => x"515473f3",
   435 => x"3873d00c",
   436 => x"7783ffe0",
   437 => x"800c02a0",
   438 => x"050d0402",
   439 => x"f4050d74",
   440 => x"70882a83",
   441 => x"fe800670",
   442 => x"72982a07",
   443 => x"72882b87",
   444 => x"fc808006",
   445 => x"73982b81",
   446 => x"f00a0671",
   447 => x"73070783",
   448 => x"ffe0800c",
   449 => x"56515351",
   450 => x"028c050d",
   451 => x"0402f805",
   452 => x"0d028e05",
   453 => x"84808080",
   454 => x"b02d7488",
   455 => x"2b077083",
   456 => x"ffff0683",
   457 => x"ffe0800c",
   458 => x"51028805",
   459 => x"0d0402f8",
   460 => x"050d7370",
   461 => x"902b7190",
   462 => x"2a0783ff",
   463 => x"e0800c52",
   464 => x"0288050d",
   465 => x"0402ec05",
   466 => x"0d800bfc",
   467 => x"800c8480",
   468 => x"80a39051",
   469 => x"84808084",
   470 => x"d62d8480",
   471 => x"808aef2d",
   472 => x"83ffe080",
   473 => x"08802e82",
   474 => x"86388480",
   475 => x"80a3a851",
   476 => x"84808084",
   477 => x"d62d8480",
   478 => x"8091d32d",
   479 => x"83ffe1a0",
   480 => x"52848080",
   481 => x"a3c05184",
   482 => x"80809ed4",
   483 => x"2d83ffe0",
   484 => x"8008802e",
   485 => x"81cd3883",
   486 => x"ffe1a00b",
   487 => x"848080a3",
   488 => x"cc525484",
   489 => x"808084d6",
   490 => x"2d805573",
   491 => x"70810555",
   492 => x"84808080",
   493 => x"b02d5372",
   494 => x"a02e80e6",
   495 => x"3872c00c",
   496 => x"72a32e81",
   497 => x"84387280",
   498 => x"c72e0981",
   499 => x"068d3884",
   500 => x"8080808c",
   501 => x"2d848080",
   502 => x"8ffd0472",
   503 => x"8a2e0981",
   504 => x"068d3884",
   505 => x"80808095",
   506 => x"2d848080",
   507 => x"8ffd0472",
   508 => x"80cc2e09",
   509 => x"81068638",
   510 => x"83ffe1a0",
   511 => x"547281df",
   512 => x"06f00570",
   513 => x"81ff0651",
   514 => x"53b87327",
   515 => x"8938ef13",
   516 => x"7081ff06",
   517 => x"51537484",
   518 => x"2b730755",
   519 => x"8480808f",
   520 => x"ab0472a3",
   521 => x"2ea33873",
   522 => x"70810555",
   523 => x"84808080",
   524 => x"b02d5372",
   525 => x"a02ef038",
   526 => x"ff147553",
   527 => x"70525484",
   528 => x"80809ed4",
   529 => x"2d74fc80",
   530 => x"0c737081",
   531 => x"05558480",
   532 => x"8080b02d",
   533 => x"53728a2e",
   534 => x"098106ed",
   535 => x"38848080",
   536 => x"8fa90484",
   537 => x"8080a3e0",
   538 => x"51848080",
   539 => x"84d62d84",
   540 => x"8080a3fc",
   541 => x"51848080",
   542 => x"84d62d80",
   543 => x"0b83ffe0",
   544 => x"800c0294",
   545 => x"050d0402",
   546 => x"e8050d77",
   547 => x"797b5855",
   548 => x"55805372",
   549 => x"7625af38",
   550 => x"74708105",
   551 => x"56848080",
   552 => x"80b02d74",
   553 => x"70810556",
   554 => x"84808080",
   555 => x"b02d5252",
   556 => x"71712e89",
   557 => x"38815184",
   558 => x"808091c8",
   559 => x"04811353",
   560 => x"84808091",
   561 => x"93048051",
   562 => x"7083ffe0",
   563 => x"800c0298",
   564 => x"050d0402",
   565 => x"d8050dff",
   566 => x"0b83fff5",
   567 => x"cc0c800b",
   568 => x"83fff5e0",
   569 => x"0c848080",
   570 => x"a4885184",
   571 => x"808084d6",
   572 => x"2d83fff1",
   573 => x"b8528051",
   574 => x"8480808c",
   575 => x"9e2d83ff",
   576 => x"e0800854",
   577 => x"83ffe080",
   578 => x"08953884",
   579 => x"8080a498",
   580 => x"51848080",
   581 => x"84d62d73",
   582 => x"55848080",
   583 => x"9a890484",
   584 => x"8080a4ac",
   585 => x"51848080",
   586 => x"84d62d80",
   587 => x"56810b83",
   588 => x"fff1ac0c",
   589 => x"88538480",
   590 => x"80a4c452",
   591 => x"83fff1ee",
   592 => x"51848080",
   593 => x"91872d83",
   594 => x"ffe08008",
   595 => x"762e0981",
   596 => x"068b3883",
   597 => x"ffe08008",
   598 => x"83fff1ac",
   599 => x"0c885384",
   600 => x"8080a4d0",
   601 => x"5283fff2",
   602 => x"8a518480",
   603 => x"8091872d",
   604 => x"83ffe080",
   605 => x"088b3883",
   606 => x"ffe08008",
   607 => x"83fff1ac",
   608 => x"0c83fff1",
   609 => x"ac085284",
   610 => x"8080a4dc",
   611 => x"51848080",
   612 => x"81f42d83",
   613 => x"fff1ac08",
   614 => x"802e81cb",
   615 => x"3883fff4",
   616 => x"fe0b8480",
   617 => x"8080b02d",
   618 => x"83fff4ff",
   619 => x"0b848080",
   620 => x"80b02d71",
   621 => x"982b7190",
   622 => x"2b0783ff",
   623 => x"f5800b84",
   624 => x"808080b0",
   625 => x"2d70882b",
   626 => x"720783ff",
   627 => x"f5810b84",
   628 => x"808080b0",
   629 => x"2d710783",
   630 => x"fff5b60b",
   631 => x"84808080",
   632 => x"b02d83ff",
   633 => x"f5b70b84",
   634 => x"808080b0",
   635 => x"2d71882b",
   636 => x"07535f54",
   637 => x"525a5657",
   638 => x"557381ab",
   639 => x"aa2e0981",
   640 => x"06953875",
   641 => x"51848080",
   642 => x"8ddb2d83",
   643 => x"ffe08008",
   644 => x"56848080",
   645 => x"94b00473",
   646 => x"82d4d52e",
   647 => x"93388480",
   648 => x"80a4f051",
   649 => x"84808084",
   650 => x"d62d8480",
   651 => x"8096bc04",
   652 => x"75528480",
   653 => x"80a59051",
   654 => x"84808081",
   655 => x"f42d83ff",
   656 => x"f1b85275",
   657 => x"51848080",
   658 => x"8c9e2d83",
   659 => x"ffe08008",
   660 => x"5583ffe0",
   661 => x"8008802e",
   662 => x"85af3884",
   663 => x"8080a5a8",
   664 => x"51848080",
   665 => x"84d62d84",
   666 => x"8080a5d0",
   667 => x"51848080",
   668 => x"81f42d88",
   669 => x"53848080",
   670 => x"a4d05283",
   671 => x"fff28a51",
   672 => x"84808091",
   673 => x"872d83ff",
   674 => x"e080088e",
   675 => x"38810b83",
   676 => x"fff5e00c",
   677 => x"84808095",
   678 => x"c8048853",
   679 => x"848080a4",
   680 => x"c45283ff",
   681 => x"f1ee5184",
   682 => x"80809187",
   683 => x"2d83ffe0",
   684 => x"8008802e",
   685 => x"93388480",
   686 => x"80a5e851",
   687 => x"84808081",
   688 => x"f42d8480",
   689 => x"8096bc04",
   690 => x"83fff5b6",
   691 => x"0b848080",
   692 => x"80b02d54",
   693 => x"7380d52e",
   694 => x"09810680",
   695 => x"df3883ff",
   696 => x"f5b70b84",
   697 => x"808080b0",
   698 => x"2d547381",
   699 => x"aa2e0981",
   700 => x"0680c938",
   701 => x"800b83ff",
   702 => x"f1b80b84",
   703 => x"808080b0",
   704 => x"2d565474",
   705 => x"81e92e83",
   706 => x"38815474",
   707 => x"81eb2e8c",
   708 => x"38805573",
   709 => x"752e0981",
   710 => x"0683ee38",
   711 => x"83fff1c3",
   712 => x"0b848080",
   713 => x"80b02d59",
   714 => x"78923883",
   715 => x"fff1c40b",
   716 => x"84808080",
   717 => x"b02d5473",
   718 => x"822e8938",
   719 => x"80558480",
   720 => x"809a8904",
   721 => x"83fff1c5",
   722 => x"0b848080",
   723 => x"80b02d70",
   724 => x"83fff5e8",
   725 => x"0cff1170",
   726 => x"83fff5dc",
   727 => x"0c545284",
   728 => x"8080a688",
   729 => x"51848080",
   730 => x"81f42d83",
   731 => x"fff1c60b",
   732 => x"84808080",
   733 => x"b02d83ff",
   734 => x"f1c70b84",
   735 => x"808080b0",
   736 => x"2d567605",
   737 => x"75828029",
   738 => x"057083ff",
   739 => x"f5d00c83",
   740 => x"fff1c80b",
   741 => x"84808080",
   742 => x"b02d7083",
   743 => x"fff5c80c",
   744 => x"83fff5e0",
   745 => x"08595758",
   746 => x"76802e81",
   747 => x"ec388853",
   748 => x"848080a4",
   749 => x"d05283ff",
   750 => x"f28a5184",
   751 => x"80809187",
   752 => x"2d785583",
   753 => x"ffe08008",
   754 => x"82bf3883",
   755 => x"fff5e808",
   756 => x"70842b83",
   757 => x"fff5b80c",
   758 => x"7083fff5",
   759 => x"e40c83ff",
   760 => x"f1dd0b84",
   761 => x"808080b0",
   762 => x"2d83fff1",
   763 => x"dc0b8480",
   764 => x"8080b02d",
   765 => x"71828029",
   766 => x"0583fff1",
   767 => x"de0b8480",
   768 => x"8080b02d",
   769 => x"70848080",
   770 => x"291283ff",
   771 => x"f1df0b84",
   772 => x"808080b0",
   773 => x"2d708180",
   774 => x"0a291270",
   775 => x"83fff1b0",
   776 => x"0c83fff5",
   777 => x"c8087129",
   778 => x"83fff5d0",
   779 => x"08057083",
   780 => x"fff5f00c",
   781 => x"83fff1e5",
   782 => x"0b848080",
   783 => x"80b02d83",
   784 => x"fff1e40b",
   785 => x"84808080",
   786 => x"b02d7182",
   787 => x"80290583",
   788 => x"fff1e60b",
   789 => x"84808080",
   790 => x"b02d7084",
   791 => x"80802912",
   792 => x"83fff1e7",
   793 => x"0b848080",
   794 => x"80b02d70",
   795 => x"982b81f0",
   796 => x"0a067205",
   797 => x"7083fff1",
   798 => x"b40cfe11",
   799 => x"7e297705",
   800 => x"83fff5d8",
   801 => x"0c525752",
   802 => x"575d5751",
   803 => x"525f525c",
   804 => x"57575784",
   805 => x"80809a87",
   806 => x"0483fff1",
   807 => x"ca0b8480",
   808 => x"8080b02d",
   809 => x"83fff1c9",
   810 => x"0b848080",
   811 => x"80b02d71",
   812 => x"82802905",
   813 => x"7083fff5",
   814 => x"b80c70a0",
   815 => x"2983ff05",
   816 => x"70892a70",
   817 => x"83fff5e4",
   818 => x"0c83fff1",
   819 => x"cf0b8480",
   820 => x"8080b02d",
   821 => x"83fff1ce",
   822 => x"0b848080",
   823 => x"80b02d71",
   824 => x"82802905",
   825 => x"7083fff1",
   826 => x"b00c7b71",
   827 => x"291e7083",
   828 => x"fff5d80c",
   829 => x"7d83fff1",
   830 => x"b40c7305",
   831 => x"83fff5f0",
   832 => x"0c555e51",
   833 => x"51555581",
   834 => x"557483ff",
   835 => x"e0800c02",
   836 => x"a8050d04",
   837 => x"02ec050d",
   838 => x"7670872c",
   839 => x"7180ff06",
   840 => x"57555383",
   841 => x"fff5e008",
   842 => x"8a387288",
   843 => x"2c7381ff",
   844 => x"06565473",
   845 => x"83fff5cc",
   846 => x"082ebc38",
   847 => x"83fff5d0",
   848 => x"08145284",
   849 => x"8080a6ac",
   850 => x"51848080",
   851 => x"81f42d83",
   852 => x"fff1b852",
   853 => x"83fff5d0",
   854 => x"08145184",
   855 => x"80808c9e",
   856 => x"2d83ffe0",
   857 => x"80085383",
   858 => x"ffe08008",
   859 => x"802e80cf",
   860 => x"387383ff",
   861 => x"f5cc0c83",
   862 => x"fff5e008",
   863 => x"802ea238",
   864 => x"74842983",
   865 => x"fff1b805",
   866 => x"70085253",
   867 => x"8480808d",
   868 => x"db2d83ff",
   869 => x"e08008f0",
   870 => x"0a065584",
   871 => x"80809bbd",
   872 => x"04741083",
   873 => x"fff1b805",
   874 => x"70848080",
   875 => x"809b2d52",
   876 => x"53848080",
   877 => x"8e8d2d83",
   878 => x"ffe08008",
   879 => x"55745372",
   880 => x"83ffe080",
   881 => x"0c029405",
   882 => x"0d0402c8",
   883 => x"050d7f61",
   884 => x"5f5c8057",
   885 => x"ff0b83ff",
   886 => x"f5cc0c83",
   887 => x"fff1b408",
   888 => x"83fff5d8",
   889 => x"08575883",
   890 => x"fff5e008",
   891 => x"772e8f38",
   892 => x"83fff5e8",
   893 => x"08842b59",
   894 => x"8480809c",
   895 => x"860483ff",
   896 => x"f5e40884",
   897 => x"2b59805a",
   898 => x"79792781",
   899 => x"ea38798f",
   900 => x"06a01858",
   901 => x"5473a438",
   902 => x"75528480",
   903 => x"80a6cc51",
   904 => x"84808081",
   905 => x"f42d83ff",
   906 => x"f1b85275",
   907 => x"51811656",
   908 => x"8480808c",
   909 => x"9e2d83ff",
   910 => x"f1b85780",
   911 => x"77848080",
   912 => x"80b02d56",
   913 => x"5474742e",
   914 => x"83388154",
   915 => x"7481e52e",
   916 => x"819c3881",
   917 => x"70750655",
   918 => x"5d73802e",
   919 => x"8190388b",
   920 => x"17848080",
   921 => x"80b02d98",
   922 => x"065b7a81",
   923 => x"81388b53",
   924 => x"7d527651",
   925 => x"84808091",
   926 => x"872d83ff",
   927 => x"e0800880",
   928 => x"ed389c17",
   929 => x"08518480",
   930 => x"808ddb2d",
   931 => x"83ffe080",
   932 => x"08841d0c",
   933 => x"9a178480",
   934 => x"80809b2d",
   935 => x"51848080",
   936 => x"8e8d2d83",
   937 => x"ffe08008",
   938 => x"83ffe080",
   939 => x"08881e0c",
   940 => x"83ffe080",
   941 => x"08555583",
   942 => x"fff5e008",
   943 => x"802ea038",
   944 => x"94178480",
   945 => x"80809b2d",
   946 => x"51848080",
   947 => x"8e8d2d83",
   948 => x"ffe08008",
   949 => x"902b83ff",
   950 => x"f00a0670",
   951 => x"16515473",
   952 => x"881d0c7a",
   953 => x"7c0c7c54",
   954 => x"8480809e",
   955 => x"c904811a",
   956 => x"5a848080",
   957 => x"9c880483",
   958 => x"fff5e008",
   959 => x"802e80c7",
   960 => x"38775184",
   961 => x"80809a94",
   962 => x"2d83ffe0",
   963 => x"800883ff",
   964 => x"e0800853",
   965 => x"848080a6",
   966 => x"ec525884",
   967 => x"808081f4",
   968 => x"2d7780ff",
   969 => x"fffff806",
   970 => x"547380ff",
   971 => x"fffff82e",
   972 => x"9638fe18",
   973 => x"83fff5e8",
   974 => x"082983ff",
   975 => x"f5f00805",
   976 => x"56848080",
   977 => x"9c860480",
   978 => x"547383ff",
   979 => x"e0800c02",
   980 => x"b8050d04",
   981 => x"02d4050d",
   982 => x"7c7e7154",
   983 => x"83fff5bc",
   984 => x"535a5784",
   985 => x"80809bca",
   986 => x"2d83ffe0",
   987 => x"800881ff",
   988 => x"06567580",
   989 => x"2e81b938",
   990 => x"848080a7",
   991 => x"84518480",
   992 => x"8084d62d",
   993 => x"83fff5c0",
   994 => x"0883ff05",
   995 => x"892a5b80",
   996 => x"70595a79",
   997 => x"7b2581b8",
   998 => x"3883fff5",
   999 => x"c408fe11",
  1000 => x"83fff5e8",
  1001 => x"082983ff",
  1002 => x"f5f00811",
  1003 => x"7a83fff5",
  1004 => x"dc080605",
  1005 => x"7a585157",
  1006 => x"5483fff5",
  1007 => x"f0085375",
  1008 => x"52848080",
  1009 => x"a7a05184",
  1010 => x"808081f4",
  1011 => x"2d785275",
  1012 => x"51848080",
  1013 => x"8c9e2d83",
  1014 => x"ffe08008",
  1015 => x"802e80e4",
  1016 => x"38848080",
  1017 => x"a7c45184",
  1018 => x"808084d6",
  1019 => x"2d811870",
  1020 => x"83fff5dc",
  1021 => x"08065758",
  1022 => x"75a33884",
  1023 => x"8080a7d4",
  1024 => x"51848080",
  1025 => x"84d62d83",
  1026 => x"fff5c408",
  1027 => x"51848080",
  1028 => x"9a942d83",
  1029 => x"ffe08008",
  1030 => x"83fff5c4",
  1031 => x"0c848019",
  1032 => x"811b5b59",
  1033 => x"7a7a24fe",
  1034 => x"f0388480",
  1035 => x"80a0d004",
  1036 => x"76528480",
  1037 => x"80a7ec51",
  1038 => x"84808081",
  1039 => x"f42d8480",
  1040 => x"80a0d204",
  1041 => x"83ffe080",
  1042 => x"08568480",
  1043 => x"80a0d204",
  1044 => x"81567583",
  1045 => x"ffe0800c",
  1046 => x"02ac050d",
  1047 => x"0483ffe0",
  1048 => x"8c080283",
  1049 => x"ffe08c0c",
  1050 => x"ff3d0d80",
  1051 => x"0b83ffe0",
  1052 => x"8c08fc05",
  1053 => x"0c83ffe0",
  1054 => x"8c088805",
  1055 => x"088106ff",
  1056 => x"11700970",
  1057 => x"83ffe08c",
  1058 => x"088c0508",
  1059 => x"0683ffe0",
  1060 => x"8c08fc05",
  1061 => x"081183ff",
  1062 => x"e08c08fc",
  1063 => x"050c83ff",
  1064 => x"e08c0888",
  1065 => x"0508812a",
  1066 => x"83ffe08c",
  1067 => x"0888050c",
  1068 => x"83ffe08c",
  1069 => x"088c0508",
  1070 => x"1083ffe0",
  1071 => x"8c088c05",
  1072 => x"0c515151",
  1073 => x"5183ffe0",
  1074 => x"8c088805",
  1075 => x"08802e84",
  1076 => x"38ffa239",
  1077 => x"83ffe08c",
  1078 => x"08fc0508",
  1079 => x"7083ffe0",
  1080 => x"800c5183",
  1081 => x"3d0d83ff",
  1082 => x"e08c0c04",
  1083 => x"00ffffff",
  1084 => x"ff00ffff",
  1085 => x"ffff00ff",
  1086 => x"ffffff00",
  1087 => x"436d645f",
  1088 => x"696e6974",
  1089 => x"0a000000",
  1090 => x"636d645f",
  1091 => x"434d4438",
  1092 => x"20726573",
  1093 => x"706f6e73",
  1094 => x"653a2025",
  1095 => x"640a0000",
  1096 => x"434d4438",
  1097 => x"5f342072",
  1098 => x"6573706f",
  1099 => x"6e73653a",
  1100 => x"2025640a",
  1101 => x"00000000",
  1102 => x"53444843",
  1103 => x"20496e69",
  1104 => x"7469616c",
  1105 => x"697a6174",
  1106 => x"696f6e20",
  1107 => x"6572726f",
  1108 => x"72210a00",
  1109 => x"434d4435",
  1110 => x"38202564",
  1111 => x"0a202000",
  1112 => x"434d4435",
  1113 => x"385f3220",
  1114 => x"25640a20",
  1115 => x"20000000",
  1116 => x"52656164",
  1117 => x"20636f6d",
  1118 => x"6d616e64",
  1119 => x"20666169",
  1120 => x"6c656420",
  1121 => x"61742025",
  1122 => x"64202825",
  1123 => x"64290a00",
  1124 => x"496e6974",
  1125 => x"69616c69",
  1126 => x"7a696e67",
  1127 => x"20534420",
  1128 => x"63617264",
  1129 => x"0a000000",
  1130 => x"48756e74",
  1131 => x"696e6720",
  1132 => x"666f7220",
  1133 => x"70617274",
  1134 => x"6974696f",
  1135 => x"6e0a0000",
  1136 => x"4d414e49",
  1137 => x"46455354",
  1138 => x"4d535400",
  1139 => x"50617273",
  1140 => x"696e6720",
  1141 => x"6d616e69",
  1142 => x"66657374",
  1143 => x"0a000000",
  1144 => x"4c6f6164",
  1145 => x"696e6720",
  1146 => x"6d616e69",
  1147 => x"66657374",
  1148 => x"20666169",
  1149 => x"6c65640a",
  1150 => x"00000000",
  1151 => x"52657475",
  1152 => x"726e696e",
  1153 => x"670a0000",
  1154 => x"52656164",
  1155 => x"696e6720",
  1156 => x"4d42520a",
  1157 => x"00000000",
  1158 => x"52656164",
  1159 => x"206f6620",
  1160 => x"4d425220",
  1161 => x"6661696c",
  1162 => x"65640a00",
  1163 => x"4d425220",
  1164 => x"73756363",
  1165 => x"65737366",
  1166 => x"756c6c79",
  1167 => x"20726561",
  1168 => x"640a0000",
  1169 => x"46415431",
  1170 => x"36202020",
  1171 => x"00000000",
  1172 => x"46415433",
  1173 => x"32202020",
  1174 => x"00000000",
  1175 => x"50617274",
  1176 => x"6974696f",
  1177 => x"6e636f75",
  1178 => x"6e742025",
  1179 => x"640a0000",
  1180 => x"4e6f2070",
  1181 => x"61727469",
  1182 => x"74696f6e",
  1183 => x"20736967",
  1184 => x"6e617475",
  1185 => x"72652066",
  1186 => x"6f756e64",
  1187 => x"0a000000",
  1188 => x"52656164",
  1189 => x"696e6720",
  1190 => x"626f6f74",
  1191 => x"20736563",
  1192 => x"746f7220",
  1193 => x"25640a00",
  1194 => x"52656164",
  1195 => x"20626f6f",
  1196 => x"74207365",
  1197 => x"63746f72",
  1198 => x"2066726f",
  1199 => x"6d206669",
  1200 => x"72737420",
  1201 => x"70617274",
  1202 => x"6974696f",
  1203 => x"6e0a0000",
  1204 => x"48756e74",
  1205 => x"696e6720",
  1206 => x"666f7220",
  1207 => x"66696c65",
  1208 => x"73797374",
  1209 => x"656d0a00",
  1210 => x"556e7375",
  1211 => x"70706f72",
  1212 => x"74656420",
  1213 => x"70617274",
  1214 => x"6974696f",
  1215 => x"6e207479",
  1216 => x"7065210d",
  1217 => x"00000000",
  1218 => x"436c7573",
  1219 => x"74657220",
  1220 => x"73697a65",
  1221 => x"3a202564",
  1222 => x"2c20436c",
  1223 => x"75737465",
  1224 => x"72206d61",
  1225 => x"736b2c20",
  1226 => x"25640a00",
  1227 => x"47657443",
  1228 => x"6c757374",
  1229 => x"65722072",
  1230 => x"65616469",
  1231 => x"6e672073",
  1232 => x"6563746f",
  1233 => x"72202564",
  1234 => x"0a000000",
  1235 => x"52656164",
  1236 => x"696e6720",
  1237 => x"64697265",
  1238 => x"63746f72",
  1239 => x"79207365",
  1240 => x"63746f72",
  1241 => x"2025640a",
  1242 => x"00000000",
  1243 => x"47657446",
  1244 => x"41544c69",
  1245 => x"6e6b2072",
  1246 => x"65747572",
  1247 => x"6e656420",
  1248 => x"25640a00",
  1249 => x"4f70656e",
  1250 => x"65642066",
  1251 => x"696c652c",
  1252 => x"206c6f61",
  1253 => x"64696e67",
  1254 => x"2e2e2e0a",
  1255 => x"00000000",
  1256 => x"52656164",
  1257 => x"696e6720",
  1258 => x"626c6f63",
  1259 => x"6b202564",
  1260 => x"20282564",
  1261 => x"2c202564",
  1262 => x"2c202564",
  1263 => x"292e2e2e",
  1264 => x"00000000",
  1265 => x"626c6f63",
  1266 => x"6b207265",
  1267 => x"61642e0a",
  1268 => x"00000000",
  1269 => x"47657474",
  1270 => x"696e6720",
  1271 => x"6e657874",
  1272 => x"20636c75",
  1273 => x"73746572",
  1274 => x"2e0a0000",
  1275 => x"43616e27",
  1276 => x"74206f70",
  1277 => x"656e2025",
  1278 => x"730a0000",
	others => x"00000000"
);

begin

process (clk)
begin
	if (clk'event and clk = '1') then
		if (from_zpu.memAWriteEnable = '1') and (from_zpu.memBWriteEnable = '1') and (from_zpu.memAAddr=from_zpu.memBAddr) and (from_zpu.memAWrite/=from_zpu.memBWrite) then
			report "write collision" severity failure;
		end if;
	
		if (from_zpu.memAWriteEnable = '1') then
			ram(to_integer(unsigned(from_zpu.memAAddr(maxAddrBitBRAM downto 2)))) := from_zpu.memAWrite;
			to_zpu.memARead <= from_zpu.memAWrite;
		else
			to_zpu.memARead <= ram(to_integer(unsigned(from_zpu.memAAddr(maxAddrBitBRAM downto 2))));
		end if;
	end if;
end process;

process (clk)
begin
	if (clk'event and clk = '1') then
		if (from_zpu.memBWriteEnable = '1') then
			ram(to_integer(unsigned(from_zpu.memBAddr(maxAddrBitBRAM downto 2)))) := from_zpu.memBWrite;
			to_zpu.memBRead <= from_zpu.memBWrite;
		else
			to_zpu.memBRead <= ram(to_integer(unsigned(from_zpu.memBAddr(maxAddrBitBRAM downto 2))));
		end if;
	end if;
end process;


end arch;

