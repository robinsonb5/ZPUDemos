-- ZPU
--
-- Copyright 2004-2008 oharboe - �yvind Harboe - oyvind.harboe@zylin.com
-- Modified by Alastair M. Robinson for the ZPUFlex project.
--
-- The FreeBSD license
-- 
-- Redistribution and use in source and binary forms, with or without
-- modification, are permitted provided that the following conditions
-- are met:
-- 
-- 1. Redistributions of source code must retain the above copyright
--    notice, this list of conditions and the following disclaimer.
-- 2. Redistributions in binary form must reproduce the above
--    copyright notice, this list of conditions and the following
--    disclaimer in the documentation and/or other materials
--    provided with the distribution.
-- 
-- THIS SOFTWARE IS PROVIDED BY THE ZPU PROJECT ``AS IS'' AND ANY
-- EXPRESS OR IMPLIED WARRANTIES, INCLUDING, BUT NOT LIMITED TO,
-- THE IMPLIED WARRANTIES OF MERCHANTABILITY AND FITNESS FOR A
-- PARTICULAR PURPOSE ARE DISCLAIMED. IN NO EVENT SHALL THE
-- ZPU PROJECT OR CONTRIBUTORS BE LIABLE FOR ANY DIRECT,
-- INDIRECT, INCIDENTAL, SPECIAL, EXEMPLARY, OR CONSEQUENTIAL DAMAGES
-- (INCLUDING, BUT NOT LIMITED TO, PROCUREMENT OF SUBSTITUTE GOODS
-- OR SERVICES; LOSS OF USE, DATA, OR PROFITS; OR BUSINESS INTERRUPTION)
-- HOWEVER CAUSED AND ON ANY THEORY OF LIABILITY, WHETHER IN CONTRACT,
-- STRICT LIABILITY, OR TORT (INCLUDING NEGLIGENCE OR OTHERWISE)
-- ARISING IN ANY WAY OUT OF THE USE OF THIS SOFTWARE, EVEN IF
-- ADVISED OF THE POSSIBILITY OF SUCH DAMAGE.
-- 
-- The views and conclusions contained in the software and documentation
-- are those of the authors and should not be interpreted as representing
-- official policies, either expressed or implied, of the ZPU Project.

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;


library work;
use work.zpu_config.all;
use work.zpupkg.all;

entity SDBootstrap_ROM is
generic
	(
		maxAddrBit : integer := maxAddrBitBRAMLimit -- Specify your actual ROM size to save LEs and unnecessary block RAM usage.
	);
port (
	clk : in std_logic;
	areset : in std_logic := '0';
	from_zpu : in ZPU_ToROM;
	to_zpu : out ZPU_FromROM
);
end SDBootstrap_ROM;

architecture arch of SDBootstrap_ROM is

type ram_type is array(natural range 0 to ((2**(maxAddrBit+1))/4)-1) of std_logic_vector(wordSize-1 downto 0);

shared variable ram : ram_type :=
(
     0 => x"0ba08080",
     1 => x"e2040000",
     2 => x"8004a080",
     3 => x"808a0471",
     4 => x"fd060872",
     5 => x"83060981",
     6 => x"05820583",
     7 => x"2b2a83ff",
     8 => x"ff065204",
     9 => x"71fc0608",
    10 => x"72830609",
    11 => x"81058305",
    12 => x"1010102a",
    13 => x"81ff0652",
    14 => x"0471fc06",
    15 => x"080ba080",
    16 => x"9ed47383",
    17 => x"06101005",
    18 => x"08067381",
    19 => x"ff067383",
    20 => x"06098105",
    21 => x"83051010",
    22 => x"102b0772",
    23 => x"fc060c51",
    24 => x"5104a080",
    25 => x"808a0ba0",
    26 => x"808d8704",
    27 => x"0002c405",
    28 => x"0d0280c0",
    29 => x"0583ffe0",
    30 => x"e05b5680",
    31 => x"76708405",
    32 => x"5808715e",
    33 => x"5e577c70",
    34 => x"84055e08",
    35 => x"58805b77",
    36 => x"982a7888",
    37 => x"2b595372",
    38 => x"8838765e",
    39 => x"a0808396",
    40 => x"047b802e",
    41 => x"81ca3880",
    42 => x"5c7280e4",
    43 => x"2e9f3872",
    44 => x"80e4268d",
    45 => x"387280e3",
    46 => x"2e80ee38",
    47 => x"a08082b6",
    48 => x"047280f3",
    49 => x"2e80cc38",
    50 => x"a08082b6",
    51 => x"04758417",
    52 => x"71087e5c",
    53 => x"56575287",
    54 => x"55739c2a",
    55 => x"74842b55",
    56 => x"5271802e",
    57 => x"83388159",
    58 => x"89722589",
    59 => x"38b71252",
    60 => x"a08081f8",
    61 => x"04b01252",
    62 => x"78802e88",
    63 => x"387151a0",
    64 => x"8083a12d",
    65 => x"ff155574",
    66 => x"8025ce38",
    67 => x"8054a080",
    68 => x"82cc0475",
    69 => x"84177108",
    70 => x"70545c57",
    71 => x"52a08083",
    72 => x"c52d7b54",
    73 => x"a08082cc",
    74 => x"04758417",
    75 => x"71085557",
    76 => x"52a08082",
    77 => x"ff04a551",
    78 => x"a08083a1",
    79 => x"2d7251a0",
    80 => x"8083a12d",
    81 => x"821757a0",
    82 => x"80838904",
    83 => x"73ff1555",
    84 => x"52807225",
    85 => x"b4387970",
    86 => x"81055ba0",
    87 => x"8080a42d",
    88 => x"705253a0",
    89 => x"8083a12d",
    90 => x"811757a0",
    91 => x"8082cc04",
    92 => x"72a52e09",
    93 => x"81068838",
    94 => x"815ca080",
    95 => x"83890472",
    96 => x"51a08083",
    97 => x"a12d8117",
    98 => x"57811b5b",
    99 => x"837b25fd",
   100 => x"fe3872fd",
   101 => x"f1387d83",
   102 => x"ffe0800c",
   103 => x"02bc050d",
   104 => x"0402f805",
   105 => x"0d7352c0",
   106 => x"0870882a",
   107 => x"70810651",
   108 => x"51517080",
   109 => x"2ef13871",
   110 => x"c00c7183",
   111 => x"ffe0800c",
   112 => x"0288050d",
   113 => x"0402e805",
   114 => x"0d775574",
   115 => x"70840556",
   116 => x"08538054",
   117 => x"72982a73",
   118 => x"882b5452",
   119 => x"71802ea2",
   120 => x"38c00870",
   121 => x"882a7081",
   122 => x"06515151",
   123 => x"70802ef1",
   124 => x"3871c00c",
   125 => x"81168115",
   126 => x"55568374",
   127 => x"25d63871",
   128 => x"ca387583",
   129 => x"ffe0800c",
   130 => x"0298050d",
   131 => x"0402f405",
   132 => x"0d747671",
   133 => x"81ff06d4",
   134 => x"0c535383",
   135 => x"fff1a008",
   136 => x"85387189",
   137 => x"2b527198",
   138 => x"2ad40c71",
   139 => x"902a7081",
   140 => x"ff06d40c",
   141 => x"5171882a",
   142 => x"7081ff06",
   143 => x"d40c5171",
   144 => x"81ff06d4",
   145 => x"0c72902a",
   146 => x"7081ff06",
   147 => x"d40c51d4",
   148 => x"087081ff",
   149 => x"06515182",
   150 => x"b8bf5270",
   151 => x"81ff2e09",
   152 => x"81069438",
   153 => x"81ff0bd4",
   154 => x"0cd40870",
   155 => x"81ff06ff",
   156 => x"14545151",
   157 => x"71e53870",
   158 => x"83ffe080",
   159 => x"0c028c05",
   160 => x"0d0402fc",
   161 => x"050d81c7",
   162 => x"5181ff0b",
   163 => x"d40cff11",
   164 => x"51708025",
   165 => x"f4380284",
   166 => x"050d0402",
   167 => x"f0050da0",
   168 => x"8085822d",
   169 => x"819c9f53",
   170 => x"805287fc",
   171 => x"80f751a0",
   172 => x"80848d2d",
   173 => x"83ffe080",
   174 => x"085483ff",
   175 => x"e0800881",
   176 => x"2e098106",
   177 => x"ab3881ff",
   178 => x"0bd40c82",
   179 => x"0a52849c",
   180 => x"80e951a0",
   181 => x"80848d2d",
   182 => x"83ffe080",
   183 => x"088d3881",
   184 => x"ff0bd40c",
   185 => x"7353a080",
   186 => x"85f704a0",
   187 => x"8085822d",
   188 => x"ff135372",
   189 => x"ffb23872",
   190 => x"83ffe080",
   191 => x"0c029005",
   192 => x"0d0402f4",
   193 => x"050d81ff",
   194 => x"0bd40ca0",
   195 => x"809ee451",
   196 => x"a08083c5",
   197 => x"2d935380",
   198 => x"5287fc80",
   199 => x"c151a080",
   200 => x"848d2d83",
   201 => x"ffe08008",
   202 => x"8d3881ff",
   203 => x"0bd40c81",
   204 => x"53a08086",
   205 => x"c104a080",
   206 => x"85822dff",
   207 => x"135372d7",
   208 => x"387283ff",
   209 => x"e0800c02",
   210 => x"8c050d04",
   211 => x"02f0050d",
   212 => x"a0808582",
   213 => x"2d83aa52",
   214 => x"849c80c8",
   215 => x"51a08084",
   216 => x"8d2d83ff",
   217 => x"e0800883",
   218 => x"ffe08008",
   219 => x"53a0809e",
   220 => x"f05254a0",
   221 => x"8080ed2d",
   222 => x"73812e09",
   223 => x"81069038",
   224 => x"d8087083",
   225 => x"ffff0654",
   226 => x"547283aa",
   227 => x"2ea338a0",
   228 => x"8086822d",
   229 => x"a08087aa",
   230 => x"048154a0",
   231 => x"8088df04",
   232 => x"a0809f88",
   233 => x"51a08080",
   234 => x"ed2d8054",
   235 => x"a08088df",
   236 => x"047352a0",
   237 => x"809fa451",
   238 => x"a08080ed",
   239 => x"2d81ff0b",
   240 => x"d40cb153",
   241 => x"a080859b",
   242 => x"2d83ffe0",
   243 => x"8008802e",
   244 => x"80f43880",
   245 => x"5287fc80",
   246 => x"fa51a080",
   247 => x"848d2d83",
   248 => x"ffe08008",
   249 => x"80d03883",
   250 => x"ffe08008",
   251 => x"52a0809f",
   252 => x"bc51a080",
   253 => x"80ed2d81",
   254 => x"ff0bd40c",
   255 => x"d40881ff",
   256 => x"067053a0",
   257 => x"809fc852",
   258 => x"54a08080",
   259 => x"ed2d81ff",
   260 => x"0bd40c81",
   261 => x"ff0bd40c",
   262 => x"81ff0bd4",
   263 => x"0c81ff0b",
   264 => x"d40c7386",
   265 => x"2a708106",
   266 => x"70565153",
   267 => x"72802eaf",
   268 => x"38a08087",
   269 => x"990483ff",
   270 => x"e0800852",
   271 => x"a0809fbc",
   272 => x"51a08080",
   273 => x"ed2d7282",
   274 => x"2efed538",
   275 => x"ff135372",
   276 => x"fef238a0",
   277 => x"809fd851",
   278 => x"a08083c5",
   279 => x"2d725473",
   280 => x"83ffe080",
   281 => x"0c029005",
   282 => x"0d0402f4",
   283 => x"050d810b",
   284 => x"83fff1a0",
   285 => x"0cd00870",
   286 => x"8f2a7081",
   287 => x"06515153",
   288 => x"72f33872",
   289 => x"d00ca080",
   290 => x"85822da0",
   291 => x"809ff051",
   292 => x"a08083c5",
   293 => x"2dd00870",
   294 => x"8f2a7081",
   295 => x"06515153",
   296 => x"72f33881",
   297 => x"0bd00c87",
   298 => x"53805284",
   299 => x"d480c051",
   300 => x"a080848d",
   301 => x"2d83ffe0",
   302 => x"8008812e",
   303 => x"09810687",
   304 => x"3883ffe0",
   305 => x"800853a0",
   306 => x"80a08051",
   307 => x"a08083c5",
   308 => x"2d72822e",
   309 => x"09810692",
   310 => x"38a080a0",
   311 => x"9451a080",
   312 => x"83c52d80",
   313 => x"53a0808a",
   314 => x"da04ff13",
   315 => x"5372ffb9",
   316 => x"38a080a0",
   317 => x"b451a080",
   318 => x"83c52da0",
   319 => x"8086cc2d",
   320 => x"83ffe080",
   321 => x"0883fff1",
   322 => x"a00c83ff",
   323 => x"e0800880",
   324 => x"2e8b38a0",
   325 => x"80a0d051",
   326 => x"a08083c5",
   327 => x"2da080a0",
   328 => x"e451a080",
   329 => x"83c52d81",
   330 => x"5287fc80",
   331 => x"d051a080",
   332 => x"848d2d81",
   333 => x"ff0bd40c",
   334 => x"d008708f",
   335 => x"2a708106",
   336 => x"51515372",
   337 => x"f33872d0",
   338 => x"0c81ff0b",
   339 => x"d40ca080",
   340 => x"a0f451a0",
   341 => x"8083c52d",
   342 => x"81537283",
   343 => x"ffe0800c",
   344 => x"028c050d",
   345 => x"04800b83",
   346 => x"ffe0800c",
   347 => x"0402e005",
   348 => x"0d797b57",
   349 => x"57805881",
   350 => x"ff0bd40c",
   351 => x"d008708f",
   352 => x"2a708106",
   353 => x"51515473",
   354 => x"f3388281",
   355 => x"0bd00c81",
   356 => x"ff0bd40c",
   357 => x"765287fc",
   358 => x"80d151a0",
   359 => x"80848d2d",
   360 => x"80dbc6df",
   361 => x"5583ffe0",
   362 => x"8008802e",
   363 => x"983883ff",
   364 => x"e0800853",
   365 => x"7652a080",
   366 => x"a18051a0",
   367 => x"8080ed2d",
   368 => x"a0808c91",
   369 => x"0481ff0b",
   370 => x"d40cd408",
   371 => x"7081ff06",
   372 => x"51547381",
   373 => x"fe2e0981",
   374 => x"069b3880",
   375 => x"ff55d808",
   376 => x"76708405",
   377 => x"580cff15",
   378 => x"55748025",
   379 => x"f1388158",
   380 => x"a0808bfb",
   381 => x"04ff1555",
   382 => x"74cb3881",
   383 => x"ff0bd40c",
   384 => x"d008708f",
   385 => x"2a708106",
   386 => x"51515473",
   387 => x"f33873d0",
   388 => x"0c7783ff",
   389 => x"e0800c02",
   390 => x"a0050d04",
   391 => x"02f4050d",
   392 => x"7470882a",
   393 => x"83fe8006",
   394 => x"7072982a",
   395 => x"0772882b",
   396 => x"87fc8080",
   397 => x"0673982b",
   398 => x"81f00a06",
   399 => x"71730707",
   400 => x"83ffe080",
   401 => x"0c565153",
   402 => x"51028c05",
   403 => x"0d0402f8",
   404 => x"050d028e",
   405 => x"05a08080",
   406 => x"a42d7498",
   407 => x"2b71902b",
   408 => x"0770902c",
   409 => x"83ffe080",
   410 => x"0c525202",
   411 => x"88050d04",
   412 => x"02f8050d",
   413 => x"7370902b",
   414 => x"71902a07",
   415 => x"83ffe080",
   416 => x"0c520288",
   417 => x"050d0402",
   418 => x"ec050d80",
   419 => x"0b870a0c",
   420 => x"a080a1a0",
   421 => x"51a08083",
   422 => x"c52da080",
   423 => x"88ea2d83",
   424 => x"ffe08008",
   425 => x"802e81e6",
   426 => x"38a080a1",
   427 => x"b851a080",
   428 => x"83c52da0",
   429 => x"808fec2d",
   430 => x"83ffe1a0",
   431 => x"52a080a1",
   432 => x"d051a080",
   433 => x"9bf52d83",
   434 => x"ffe08008",
   435 => x"802e81be",
   436 => x"3883ffe1",
   437 => x"a00ba080",
   438 => x"a1dc5254",
   439 => x"a08083c5",
   440 => x"2d805573",
   441 => x"70810555",
   442 => x"a08080a4",
   443 => x"2d5372a0",
   444 => x"2e80de38",
   445 => x"72a32e80",
   446 => x"fd387280",
   447 => x"c72e0981",
   448 => x"068b38a0",
   449 => x"8080882d",
   450 => x"a0808ead",
   451 => x"04728a2e",
   452 => x"0981068b",
   453 => x"38a08080",
   454 => x"8a2da080",
   455 => x"8ead0472",
   456 => x"80cc2e09",
   457 => x"81068638",
   458 => x"83ffe1a0",
   459 => x"547281df",
   460 => x"06f00570",
   461 => x"81ff0651",
   462 => x"53b87327",
   463 => x"8938ef13",
   464 => x"7081ff06",
   465 => x"51537484",
   466 => x"2b730755",
   467 => x"a0808de3",
   468 => x"0472a32e",
   469 => x"a1387370",
   470 => x"810555a0",
   471 => x"8080a42d",
   472 => x"5372a02e",
   473 => x"f138ff14",
   474 => x"75537052",
   475 => x"54a0809b",
   476 => x"f52d7487",
   477 => x"0a0c7370",
   478 => x"810555a0",
   479 => x"8080a42d",
   480 => x"53728a2e",
   481 => x"098106ee",
   482 => x"38a0808d",
   483 => x"e104a080",
   484 => x"a1f051a0",
   485 => x"8083c52d",
   486 => x"800b83ff",
   487 => x"e0800c02",
   488 => x"94050d04",
   489 => x"02e8050d",
   490 => x"77797b58",
   491 => x"55558053",
   492 => x"727625ab",
   493 => x"38747081",
   494 => x"0556a080",
   495 => x"80a42d74",
   496 => x"70810556",
   497 => x"a08080a4",
   498 => x"2d525271",
   499 => x"712e8838",
   500 => x"8151a080",
   501 => x"8fe10481",
   502 => x"1353a080",
   503 => x"8fb00480",
   504 => x"517083ff",
   505 => x"e0800c02",
   506 => x"98050d04",
   507 => x"02d8050d",
   508 => x"ff0b83ff",
   509 => x"f5cc0c80",
   510 => x"0b83fff5",
   511 => x"e00ca080",
   512 => x"a1fc51a0",
   513 => x"8083c52d",
   514 => x"83fff1b8",
   515 => x"528051a0",
   516 => x"808aed2d",
   517 => x"83ffe080",
   518 => x"085483ff",
   519 => x"e0800892",
   520 => x"38a080a2",
   521 => x"8c51a080",
   522 => x"83c52d73",
   523 => x"55a08097",
   524 => x"d004a080",
   525 => x"a2a051a0",
   526 => x"8083c52d",
   527 => x"8056810b",
   528 => x"83fff1ac",
   529 => x"0c8853a0",
   530 => x"80a2b852",
   531 => x"83fff1ee",
   532 => x"51a0808f",
   533 => x"a42d83ff",
   534 => x"e0800876",
   535 => x"2e098106",
   536 => x"8b3883ff",
   537 => x"e0800883",
   538 => x"fff1ac0c",
   539 => x"8853a080",
   540 => x"a2c45283",
   541 => x"fff28a51",
   542 => x"a0808fa4",
   543 => x"2d83ffe0",
   544 => x"80088b38",
   545 => x"83ffe080",
   546 => x"0883fff1",
   547 => x"ac0c83ff",
   548 => x"f1ac0852",
   549 => x"a080a2d0",
   550 => x"51a08080",
   551 => x"ed2d83ff",
   552 => x"f1ac0880",
   553 => x"2e81bb38",
   554 => x"83fff4fe",
   555 => x"0ba08080",
   556 => x"a42d83ff",
   557 => x"f4ff0ba0",
   558 => x"8080a42d",
   559 => x"71982b71",
   560 => x"902b0783",
   561 => x"fff5800b",
   562 => x"a08080a4",
   563 => x"2d70882b",
   564 => x"720783ff",
   565 => x"f5810ba0",
   566 => x"8080a42d",
   567 => x"710783ff",
   568 => x"f5b60ba0",
   569 => x"8080a42d",
   570 => x"83fff5b7",
   571 => x"0ba08080",
   572 => x"a42d7188",
   573 => x"2b07535f",
   574 => x"54525a56",
   575 => x"57557381",
   576 => x"abaa2e09",
   577 => x"81069338",
   578 => x"7551a080",
   579 => x"8c9c2d83",
   580 => x"ffe08008",
   581 => x"56a08092",
   582 => x"b0047382",
   583 => x"d4d52e90",
   584 => x"38a080a2",
   585 => x"e451a080",
   586 => x"83c52da0",
   587 => x"8094a804",
   588 => x"7552a080",
   589 => x"a38451a0",
   590 => x"8080ed2d",
   591 => x"83fff1b8",
   592 => x"527551a0",
   593 => x"808aed2d",
   594 => x"83ffe080",
   595 => x"085583ff",
   596 => x"e0800880",
   597 => x"2e84f938",
   598 => x"a080a39c",
   599 => x"51a08083",
   600 => x"c52da080",
   601 => x"a3c451a0",
   602 => x"8080ed2d",
   603 => x"8853a080",
   604 => x"a2c45283",
   605 => x"fff28a51",
   606 => x"a0808fa4",
   607 => x"2d83ffe0",
   608 => x"80088d38",
   609 => x"810b83ff",
   610 => x"f5e00ca0",
   611 => x"8093b904",
   612 => x"8853a080",
   613 => x"a2b85283",
   614 => x"fff1ee51",
   615 => x"a0808fa4",
   616 => x"2d83ffe0",
   617 => x"8008802e",
   618 => x"9038a080",
   619 => x"a3dc51a0",
   620 => x"8080ed2d",
   621 => x"a08094a8",
   622 => x"0483fff5",
   623 => x"b60ba080",
   624 => x"80a42d54",
   625 => x"7380d52e",
   626 => x"09810680",
   627 => x"db3883ff",
   628 => x"f5b70ba0",
   629 => x"8080a42d",
   630 => x"547381aa",
   631 => x"2e098106",
   632 => x"80c63880",
   633 => x"0b83fff1",
   634 => x"b80ba080",
   635 => x"80a42d56",
   636 => x"547481e9",
   637 => x"2e833881",
   638 => x"547481eb",
   639 => x"2e8c3880",
   640 => x"5573752e",
   641 => x"09810683",
   642 => x"c73883ff",
   643 => x"f1c30ba0",
   644 => x"8080a42d",
   645 => x"55749138",
   646 => x"83fff1c4",
   647 => x"0ba08080",
   648 => x"a42d5473",
   649 => x"822e8838",
   650 => x"8055a080",
   651 => x"97d00483",
   652 => x"fff1c50b",
   653 => x"a08080a4",
   654 => x"2d7083ff",
   655 => x"f5e80cff",
   656 => x"0583fff5",
   657 => x"dc0c83ff",
   658 => x"f1c60ba0",
   659 => x"8080a42d",
   660 => x"83fff1c7",
   661 => x"0ba08080",
   662 => x"a42d5876",
   663 => x"05778280",
   664 => x"29057083",
   665 => x"fff5d00c",
   666 => x"83fff1c8",
   667 => x"0ba08080",
   668 => x"a42d7083",
   669 => x"fff5c80c",
   670 => x"83fff5e0",
   671 => x"08595758",
   672 => x"76802e81",
   673 => x"df388853",
   674 => x"a080a2c4",
   675 => x"5283fff2",
   676 => x"8a51a080",
   677 => x"8fa42d83",
   678 => x"ffe08008",
   679 => x"82b23883",
   680 => x"fff5e808",
   681 => x"70842b83",
   682 => x"fff5b80c",
   683 => x"7083fff5",
   684 => x"e40c83ff",
   685 => x"f1dd0ba0",
   686 => x"8080a42d",
   687 => x"83fff1dc",
   688 => x"0ba08080",
   689 => x"a42d7182",
   690 => x"80290583",
   691 => x"fff1de0b",
   692 => x"a08080a4",
   693 => x"2d708480",
   694 => x"80291283",
   695 => x"fff1df0b",
   696 => x"a08080a4",
   697 => x"2d708180",
   698 => x"0a291270",
   699 => x"83fff1b0",
   700 => x"0c83fff5",
   701 => x"c8087129",
   702 => x"83fff5d0",
   703 => x"08057083",
   704 => x"fff5f00c",
   705 => x"83fff1e5",
   706 => x"0ba08080",
   707 => x"a42d83ff",
   708 => x"f1e40ba0",
   709 => x"8080a42d",
   710 => x"71828029",
   711 => x"0583fff1",
   712 => x"e60ba080",
   713 => x"80a42d70",
   714 => x"84808029",
   715 => x"1283fff1",
   716 => x"e70ba080",
   717 => x"80a42d70",
   718 => x"982b81f0",
   719 => x"0a067205",
   720 => x"7083fff1",
   721 => x"b40cfe11",
   722 => x"7e297705",
   723 => x"83fff5d8",
   724 => x"0c525952",
   725 => x"43545e51",
   726 => x"5259525d",
   727 => x"575957a0",
   728 => x"8097ce04",
   729 => x"83fff1ca",
   730 => x"0ba08080",
   731 => x"a42d83ff",
   732 => x"f1c90ba0",
   733 => x"8080a42d",
   734 => x"71828029",
   735 => x"057083ff",
   736 => x"f5b80c70",
   737 => x"a02983ff",
   738 => x"0570892a",
   739 => x"7083fff5",
   740 => x"e40c83ff",
   741 => x"f1cf0ba0",
   742 => x"8080a42d",
   743 => x"83fff1ce",
   744 => x"0ba08080",
   745 => x"a42d7182",
   746 => x"80290570",
   747 => x"83fff1b0",
   748 => x"0c7b7129",
   749 => x"1e7083ff",
   750 => x"f5d80c7d",
   751 => x"83fff1b4",
   752 => x"0c730583",
   753 => x"fff5f00c",
   754 => x"555e5151",
   755 => x"55558155",
   756 => x"7483ffe0",
   757 => x"800c02a8",
   758 => x"050d0402",
   759 => x"ec050d76",
   760 => x"70872c71",
   761 => x"80ff0657",
   762 => x"555383ff",
   763 => x"f5e0088a",
   764 => x"3872882c",
   765 => x"7381ff06",
   766 => x"56547383",
   767 => x"fff5cc08",
   768 => x"2ea83883",
   769 => x"fff1b852",
   770 => x"83fff5d0",
   771 => x"081451a0",
   772 => x"808aed2d",
   773 => x"83ffe080",
   774 => x"085383ff",
   775 => x"e0800880",
   776 => x"2e80cb38",
   777 => x"7383fff5",
   778 => x"cc0c83ff",
   779 => x"f5e00880",
   780 => x"2ea03874",
   781 => x"842983ff",
   782 => x"f1b80570",
   783 => x"085253a0",
   784 => x"808c9c2d",
   785 => x"83ffe080",
   786 => x"08f00a06",
   787 => x"55a08098",
   788 => x"ec047410",
   789 => x"83fff1b8",
   790 => x"0570a080",
   791 => x"808f2d52",
   792 => x"53a0808c",
   793 => x"ce2d83ff",
   794 => x"e0800855",
   795 => x"74537283",
   796 => x"ffe0800c",
   797 => x"0294050d",
   798 => x"0402cc05",
   799 => x"0d7e605e",
   800 => x"5b8056ff",
   801 => x"0b83fff5",
   802 => x"cc0c83ff",
   803 => x"f1b40883",
   804 => x"fff5d808",
   805 => x"565783ff",
   806 => x"f5e00876",
   807 => x"2e8e3883",
   808 => x"fff5e808",
   809 => x"842b59a0",
   810 => x"8099b404",
   811 => x"83fff5e4",
   812 => x"08842b59",
   813 => x"805a7979",
   814 => x"2781e138",
   815 => x"798f06a0",
   816 => x"17575473",
   817 => x"a1387452",
   818 => x"a080a3fc",
   819 => x"51a08080",
   820 => x"ed2d83ff",
   821 => x"f1b85274",
   822 => x"51811555",
   823 => x"a0808aed",
   824 => x"2d83fff1",
   825 => x"b8568076",
   826 => x"a08080a4",
   827 => x"2d555873",
   828 => x"782e8338",
   829 => x"81587381",
   830 => x"e52e8198",
   831 => x"38817079",
   832 => x"06555c73",
   833 => x"802e818c",
   834 => x"388b16a0",
   835 => x"8080a42d",
   836 => x"98065877",
   837 => x"80fe388b",
   838 => x"537c5275",
   839 => x"51a0808f",
   840 => x"a42d83ff",
   841 => x"e0800880",
   842 => x"eb389c16",
   843 => x"0851a080",
   844 => x"8c9c2d83",
   845 => x"ffe08008",
   846 => x"841c0c9a",
   847 => x"16a08080",
   848 => x"8f2d51a0",
   849 => x"808cce2d",
   850 => x"83ffe080",
   851 => x"0883ffe0",
   852 => x"80085555",
   853 => x"83fff5e0",
   854 => x"08802e9e",
   855 => x"389416a0",
   856 => x"80808f2d",
   857 => x"51a0808c",
   858 => x"ce2d83ff",
   859 => x"e0800890",
   860 => x"2b83fff0",
   861 => x"0a067016",
   862 => x"51547388",
   863 => x"1c0c777b",
   864 => x"0c7c52a0",
   865 => x"80a49c51",
   866 => x"a08080ed",
   867 => x"2d7b54a0",
   868 => x"809bea04",
   869 => x"811a5aa0",
   870 => x"8099b604",
   871 => x"83fff5e0",
   872 => x"08802e80",
   873 => x"c3387651",
   874 => x"a08097db",
   875 => x"2d83ffe0",
   876 => x"800883ff",
   877 => x"e0800853",
   878 => x"a080a4b0",
   879 => x"5257a080",
   880 => x"80ed2d76",
   881 => x"80ffffff",
   882 => x"f8065473",
   883 => x"80ffffff",
   884 => x"f82e9538",
   885 => x"fe1783ff",
   886 => x"f5e80829",
   887 => x"83fff5f0",
   888 => x"080555a0",
   889 => x"8099b404",
   890 => x"80547383",
   891 => x"ffe0800c",
   892 => x"02b4050d",
   893 => x"0402e405",
   894 => x"0d787a71",
   895 => x"5483fff5",
   896 => x"bc535555",
   897 => x"a08098f9",
   898 => x"2d83ffe0",
   899 => x"800881ff",
   900 => x"06537280",
   901 => x"2e818338",
   902 => x"a080a4c8",
   903 => x"51a08083",
   904 => x"c52d83ff",
   905 => x"f5c00883",
   906 => x"ff05892a",
   907 => x"57807056",
   908 => x"56757725",
   909 => x"81803883",
   910 => x"fff5c408",
   911 => x"fe0583ff",
   912 => x"f5e80829",
   913 => x"83fff5f0",
   914 => x"08117683",
   915 => x"fff5dc08",
   916 => x"06057554",
   917 => x"5253a080",
   918 => x"8aed2d83",
   919 => x"ffe08008",
   920 => x"802e80c7",
   921 => x"38811570",
   922 => x"83fff5dc",
   923 => x"08065455",
   924 => x"72963883",
   925 => x"fff5c408",
   926 => x"51a08097",
   927 => x"db2d83ff",
   928 => x"e0800883",
   929 => x"fff5c40c",
   930 => x"84801481",
   931 => x"17575476",
   932 => x"7624ffa3",
   933 => x"38a0809d",
   934 => x"b6047452",
   935 => x"a080a4e4",
   936 => x"51a08080",
   937 => x"ed2da080",
   938 => x"9db80483",
   939 => x"ffe08008",
   940 => x"53a0809d",
   941 => x"b8048153",
   942 => x"7283ffe0",
   943 => x"800c029c",
   944 => x"050d0483",
   945 => x"ffe08c08",
   946 => x"0283ffe0",
   947 => x"8c0cff3d",
   948 => x"0d800b83",
   949 => x"ffe08c08",
   950 => x"fc050c83",
   951 => x"ffe08c08",
   952 => x"88050881",
   953 => x"06ff1170",
   954 => x"097083ff",
   955 => x"e08c088c",
   956 => x"05080683",
   957 => x"ffe08c08",
   958 => x"fc050811",
   959 => x"83ffe08c",
   960 => x"08fc050c",
   961 => x"83ffe08c",
   962 => x"08880508",
   963 => x"812a83ff",
   964 => x"e08c0888",
   965 => x"050c83ff",
   966 => x"e08c088c",
   967 => x"05081083",
   968 => x"ffe08c08",
   969 => x"8c050c51",
   970 => x"51515183",
   971 => x"ffe08c08",
   972 => x"88050880",
   973 => x"2e8438ff",
   974 => x"a23983ff",
   975 => x"e08c08fc",
   976 => x"05087083",
   977 => x"ffe0800c",
   978 => x"51833d0d",
   979 => x"83ffe08c",
   980 => x"0c040000",
   981 => x"00ffffff",
   982 => x"ff00ffff",
   983 => x"ffff00ff",
   984 => x"ffffff00",
   985 => x"436d645f",
   986 => x"696e6974",
   987 => x"0a000000",
   988 => x"636d645f",
   989 => x"434d4438",
   990 => x"20726573",
   991 => x"706f6e73",
   992 => x"653a2025",
   993 => x"640a0000",
   994 => x"53444843",
   995 => x"20496e69",
   996 => x"7469616c",
   997 => x"697a6174",
   998 => x"696f6e20",
   999 => x"6572726f",
  1000 => x"72210a00",
  1001 => x"434d4438",
  1002 => x"5f342072",
  1003 => x"6573706f",
  1004 => x"6e73653a",
  1005 => x"2025640a",
  1006 => x"00000000",
  1007 => x"434d4435",
  1008 => x"38202564",
  1009 => x"0a202000",
  1010 => x"434d4435",
  1011 => x"385f3220",
  1012 => x"25640a20",
  1013 => x"20000000",
  1014 => x"44657465",
  1015 => x"726d696e",
  1016 => x"65642053",
  1017 => x"44484320",
  1018 => x"73746174",
  1019 => x"75730a00",
  1020 => x"41637469",
  1021 => x"76617469",
  1022 => x"6e672043",
  1023 => x"530a0000",
  1024 => x"53656e74",
  1025 => x"20726573",
  1026 => x"65742063",
  1027 => x"6f6d6d61",
  1028 => x"6e640a00",
  1029 => x"53442063",
  1030 => x"61726420",
  1031 => x"696e6974",
  1032 => x"69616c69",
  1033 => x"7a617469",
  1034 => x"6f6e2065",
  1035 => x"72726f72",
  1036 => x"210a0000",
  1037 => x"43617264",
  1038 => x"20726573",
  1039 => x"706f6e64",
  1040 => x"65642074",
  1041 => x"6f207265",
  1042 => x"7365740a",
  1043 => x"00000000",
  1044 => x"53444843",
  1045 => x"20636172",
  1046 => x"64206465",
  1047 => x"74656374",
  1048 => x"65640a00",
  1049 => x"53656e64",
  1050 => x"696e6720",
  1051 => x"636d6431",
  1052 => x"360a0000",
  1053 => x"496e6974",
  1054 => x"20646f6e",
  1055 => x"650a0000",
  1056 => x"52656164",
  1057 => x"20636f6d",
  1058 => x"6d616e64",
  1059 => x"20666169",
  1060 => x"6c656420",
  1061 => x"61742025",
  1062 => x"64202825",
  1063 => x"64290a00",
  1064 => x"496e6974",
  1065 => x"69616c69",
  1066 => x"7a696e67",
  1067 => x"20534420",
  1068 => x"63617264",
  1069 => x"0a000000",
  1070 => x"48756e74",
  1071 => x"696e6720",
  1072 => x"666f7220",
  1073 => x"70617274",
  1074 => x"6974696f",
  1075 => x"6e0a0000",
  1076 => x"4d414e49",
  1077 => x"46455354",
  1078 => x"4d535400",
  1079 => x"50617273",
  1080 => x"696e6720",
  1081 => x"6d616e69",
  1082 => x"66657374",
  1083 => x"0a000000",
  1084 => x"52657475",
  1085 => x"726e696e",
  1086 => x"670a0000",
  1087 => x"52656164",
  1088 => x"696e6720",
  1089 => x"4d42520a",
  1090 => x"00000000",
  1091 => x"52656164",
  1092 => x"206f6620",
  1093 => x"4d425220",
  1094 => x"6661696c",
  1095 => x"65640a00",
  1096 => x"4d425220",
  1097 => x"73756363",
  1098 => x"65737366",
  1099 => x"756c6c79",
  1100 => x"20726561",
  1101 => x"640a0000",
  1102 => x"46415431",
  1103 => x"36202020",
  1104 => x"00000000",
  1105 => x"46415433",
  1106 => x"32202020",
  1107 => x"00000000",
  1108 => x"50617274",
  1109 => x"6974696f",
  1110 => x"6e636f75",
  1111 => x"6e742025",
  1112 => x"640a0000",
  1113 => x"4e6f2070",
  1114 => x"61727469",
  1115 => x"74696f6e",
  1116 => x"20736967",
  1117 => x"6e617475",
  1118 => x"72652066",
  1119 => x"6f756e64",
  1120 => x"0a000000",
  1121 => x"52656164",
  1122 => x"696e6720",
  1123 => x"626f6f74",
  1124 => x"20736563",
  1125 => x"746f7220",
  1126 => x"25640a00",
  1127 => x"52656164",
  1128 => x"20626f6f",
  1129 => x"74207365",
  1130 => x"63746f72",
  1131 => x"2066726f",
  1132 => x"6d206669",
  1133 => x"72737420",
  1134 => x"70617274",
  1135 => x"6974696f",
  1136 => x"6e0a0000",
  1137 => x"48756e74",
  1138 => x"696e6720",
  1139 => x"666f7220",
  1140 => x"66696c65",
  1141 => x"73797374",
  1142 => x"656d0a00",
  1143 => x"556e7375",
  1144 => x"70706f72",
  1145 => x"74656420",
  1146 => x"70617274",
  1147 => x"6974696f",
  1148 => x"6e207479",
  1149 => x"7065210d",
  1150 => x"00000000",
  1151 => x"52656164",
  1152 => x"696e6720",
  1153 => x"64697265",
  1154 => x"63746f72",
  1155 => x"79207365",
  1156 => x"63746f72",
  1157 => x"2025640a",
  1158 => x"00000000",
  1159 => x"66696c65",
  1160 => x"20222573",
  1161 => x"2220666f",
  1162 => x"756e640d",
  1163 => x"00000000",
  1164 => x"47657446",
  1165 => x"41544c69",
  1166 => x"6e6b2072",
  1167 => x"65747572",
  1168 => x"6e656420",
  1169 => x"25640a00",
  1170 => x"4f70656e",
  1171 => x"65642066",
  1172 => x"696c652c",
  1173 => x"206c6f61",
  1174 => x"64696e67",
  1175 => x"2e2e2e0a",
  1176 => x"00000000",
  1177 => x"43616e27",
  1178 => x"74206f70",
  1179 => x"656e2025",
  1180 => x"730a0000",
	others => x"00000000"
);

begin

process (clk)
begin
	if (clk'event and clk = '1') then
		if (from_zpu.memAWriteEnable = '1') and (from_zpu.memBWriteEnable = '1') and (from_zpu.memAAddr=from_zpu.memBAddr) and (from_zpu.memAWrite/=from_zpu.memBWrite) then
			report "write collision" severity failure;
		end if;
	
		if (from_zpu.memAWriteEnable = '1') then
			ram(to_integer(unsigned(from_zpu.memAAddr(maxAddrBit downto 2)))) := from_zpu.memAWrite;
			to_zpu.memARead <= from_zpu.memAWrite;
		else
			to_zpu.memARead <= ram(to_integer(unsigned(from_zpu.memAAddr(maxAddrBit downto 2))));
		end if;
	end if;
end process;

process (clk)
begin
	if (clk'event and clk = '1') then
		if (from_zpu.memBWriteEnable = '1') then
			ram(to_integer(unsigned(from_zpu.memBAddr(maxAddrBit downto 2)))) := from_zpu.memBWrite;
			to_zpu.memBRead <= from_zpu.memBWrite;
		else
			to_zpu.memBRead <= ram(to_integer(unsigned(from_zpu.memBAddr(maxAddrBit downto 2))));
		end if;
	end if;
end process;


end arch;

