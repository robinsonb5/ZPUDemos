-- ZPU
--
-- Copyright 2004-2008 oharboe - �yvind Harboe - oyvind.harboe@zylin.com
-- Modified by Alastair M. Robinson for the ZPUFlex project.
--
-- The FreeBSD license
-- 
-- Redistribution and use in source and binary forms, with or without
-- modification, are permitted provided that the following conditions
-- are met:
-- 
-- 1. Redistributions of source code must retain the above copyright
--    notice, this list of conditions and the following disclaimer.
-- 2. Redistributions in binary form must reproduce the above
--    copyright notice, this list of conditions and the following
--    disclaimer in the documentation and/or other materials
--    provided with the distribution.
-- 
-- THIS SOFTWARE IS PROVIDED BY THE ZPU PROJECT ``AS IS'' AND ANY
-- EXPRESS OR IMPLIED WARRANTIES, INCLUDING, BUT NOT LIMITED TO,
-- THE IMPLIED WARRANTIES OF MERCHANTABILITY AND FITNESS FOR A
-- PARTICULAR PURPOSE ARE DISCLAIMED. IN NO EVENT SHALL THE
-- ZPU PROJECT OR CONTRIBUTORS BE LIABLE FOR ANY DIRECT,
-- INDIRECT, INCIDENTAL, SPECIAL, EXEMPLARY, OR CONSEQUENTIAL DAMAGES
-- (INCLUDING, BUT NOT LIMITED TO, PROCUREMENT OF SUBSTITUTE GOODS
-- OR SERVICES; LOSS OF USE, DATA, OR PROFITS; OR BUSINESS INTERRUPTION)
-- HOWEVER CAUSED AND ON ANY THEORY OF LIABILITY, WHETHER IN CONTRACT,
-- STRICT LIABILITY, OR TORT (INCLUDING NEGLIGENCE OR OTHERWISE)
-- ARISING IN ANY WAY OUT OF THE USE OF THIS SOFTWARE, EVEN IF
-- ADVISED OF THE POSSIBILITY OF SUCH DAMAGE.
-- 
-- The views and conclusions contained in the software and documentation
-- are those of the authors and should not be interpreted as representing
-- official policies, either expressed or implied, of the ZPU Project.

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;


library work;
use work.zpu_config.all;
use work.zpupkg.all;

entity Dhrystone_fast_ROM is
generic
	(
		maxAddrBit : integer := maxAddrBitBRAMLimit -- Specify your actual ROM size to save LEs and unnecessary block RAM usage.
	);
port (
	clk : in std_logic;
	areset : in std_logic := '0';
	from_zpu : in ZPU_ToROM;
	to_zpu : out ZPU_FromROM
);
end Dhrystone_fast_ROM;

architecture arch of Dhrystone_fast_ROM is

type ram_type is array(natural range 0 to ((2**(maxAddrBit+1))/4)-1) of std_logic_vector(wordSize-1 downto 0);

shared variable ram : ram_type :=
(
     0 => x"0b0b0b88",
     1 => x"dd040000",
     2 => x"00000000",
     3 => x"00000000",
     4 => x"00000000",
     5 => x"00000000",
     6 => x"00000000",
     7 => x"00000000",
     8 => x"04000000",
     9 => x"00000000",
    10 => x"00000000",
    11 => x"00000000",
    12 => x"00000000",
    13 => x"00000000",
    14 => x"00000000",
    15 => x"00000000",
    16 => x"71fd0608",
    17 => x"72830609",
    18 => x"81058205",
    19 => x"832b2a83",
    20 => x"ffff0652",
    21 => x"04000000",
    22 => x"00000000",
    23 => x"00000000",
    24 => x"71fd0608",
    25 => x"83ffff73",
    26 => x"83060981",
    27 => x"05820583",
    28 => x"2b2b0906",
    29 => x"7383ffff",
    30 => x"0b0b0b0b",
    31 => x"83a50400",
    32 => x"72098105",
    33 => x"72057373",
    34 => x"09060906",
    35 => x"73097306",
    36 => x"070a8106",
    37 => x"53510400",
    38 => x"00000000",
    39 => x"00000000",
    40 => x"72722473",
    41 => x"732e0753",
    42 => x"51040000",
    43 => x"00000000",
    44 => x"00000000",
    45 => x"00000000",
    46 => x"00000000",
    47 => x"00000000",
    48 => x"71737109",
    49 => x"71068106",
    50 => x"09810572",
    51 => x"0a100a72",
    52 => x"0a100a31",
    53 => x"050a8106",
    54 => x"51515351",
    55 => x"04000000",
    56 => x"72722673",
    57 => x"732e0753",
    58 => x"51040000",
    59 => x"00000000",
    60 => x"00000000",
    61 => x"00000000",
    62 => x"00000000",
    63 => x"00000000",
    64 => x"00000000",
    65 => x"00000000",
    66 => x"00000000",
    67 => x"00000000",
    68 => x"00000000",
    69 => x"00000000",
    70 => x"00000000",
    71 => x"00000000",
    72 => x"0b0b0b88",
    73 => x"ba040000",
    74 => x"00000000",
    75 => x"00000000",
    76 => x"00000000",
    77 => x"00000000",
    78 => x"00000000",
    79 => x"00000000",
    80 => x"720a722b",
    81 => x"0a535104",
    82 => x"00000000",
    83 => x"00000000",
    84 => x"00000000",
    85 => x"00000000",
    86 => x"00000000",
    87 => x"00000000",
    88 => x"72729f06",
    89 => x"0981050b",
    90 => x"0b0b889f",
    91 => x"05040000",
    92 => x"00000000",
    93 => x"00000000",
    94 => x"00000000",
    95 => x"00000000",
    96 => x"72722aff",
    97 => x"739f062a",
    98 => x"0974090a",
    99 => x"8106ff05",
   100 => x"06075351",
   101 => x"04000000",
   102 => x"00000000",
   103 => x"00000000",
   104 => x"71715351",
   105 => x"04067383",
   106 => x"06098105",
   107 => x"8205832b",
   108 => x"0b2b0772",
   109 => x"fc060c51",
   110 => x"51040000",
   111 => x"00000000",
   112 => x"72098105",
   113 => x"72050970",
   114 => x"81050906",
   115 => x"0a810653",
   116 => x"51040000",
   117 => x"00000000",
   118 => x"00000000",
   119 => x"00000000",
   120 => x"72098105",
   121 => x"72050970",
   122 => x"81050906",
   123 => x"0a098106",
   124 => x"53510400",
   125 => x"00000000",
   126 => x"00000000",
   127 => x"00000000",
   128 => x"71098105",
   129 => x"52040000",
   130 => x"00000000",
   131 => x"00000000",
   132 => x"00000000",
   133 => x"00000000",
   134 => x"00000000",
   135 => x"00000000",
   136 => x"72720981",
   137 => x"05055351",
   138 => x"04000000",
   139 => x"00000000",
   140 => x"00000000",
   141 => x"00000000",
   142 => x"00000000",
   143 => x"00000000",
   144 => x"72097206",
   145 => x"73730906",
   146 => x"07535104",
   147 => x"00000000",
   148 => x"00000000",
   149 => x"00000000",
   150 => x"00000000",
   151 => x"00000000",
   152 => x"71fc0608",
   153 => x"72830609",
   154 => x"81058305",
   155 => x"1010102a",
   156 => x"81ff0652",
   157 => x"04000000",
   158 => x"00000000",
   159 => x"00000000",
   160 => x"71fc0608",
   161 => x"0b0b0ba0",
   162 => x"90738306",
   163 => x"10100508",
   164 => x"060b0b0b",
   165 => x"88a20400",
   166 => x"00000000",
   167 => x"00000000",
   168 => x"88088c08",
   169 => x"90087575",
   170 => x"0b0b0b99",
   171 => x"822d5050",
   172 => x"88085690",
   173 => x"0c8c0c88",
   174 => x"0c510400",
   175 => x"00000000",
   176 => x"88088c08",
   177 => x"90087575",
   178 => x"0b0b0b9a",
   179 => x"b42d5050",
   180 => x"88085690",
   181 => x"0c8c0c88",
   182 => x"0c510400",
   183 => x"00000000",
   184 => x"72097081",
   185 => x"0509060a",
   186 => x"8106ff05",
   187 => x"70547106",
   188 => x"73097274",
   189 => x"05ff0506",
   190 => x"07515151",
   191 => x"04000000",
   192 => x"72097081",
   193 => x"0509060a",
   194 => x"098106ff",
   195 => x"05705471",
   196 => x"06730972",
   197 => x"7405ff05",
   198 => x"06075151",
   199 => x"51040000",
   200 => x"05ff0504",
   201 => x"00000000",
   202 => x"00000000",
   203 => x"00000000",
   204 => x"00000000",
   205 => x"00000000",
   206 => x"00000000",
   207 => x"00000000",
   208 => x"04000000",
   209 => x"00000000",
   210 => x"00000000",
   211 => x"00000000",
   212 => x"00000000",
   213 => x"00000000",
   214 => x"00000000",
   215 => x"00000000",
   216 => x"71810552",
   217 => x"04000000",
   218 => x"00000000",
   219 => x"00000000",
   220 => x"00000000",
   221 => x"00000000",
   222 => x"00000000",
   223 => x"00000000",
   224 => x"00000000",
   225 => x"00000000",
   226 => x"00000000",
   227 => x"00000000",
   228 => x"00000000",
   229 => x"00000000",
   230 => x"00000000",
   231 => x"00000000",
   232 => x"02840572",
   233 => x"10100552",
   234 => x"04000000",
   235 => x"00000000",
   236 => x"00000000",
   237 => x"00000000",
   238 => x"00000000",
   239 => x"00000000",
   240 => x"00000000",
   241 => x"00000000",
   242 => x"00000000",
   243 => x"00000000",
   244 => x"00000000",
   245 => x"00000000",
   246 => x"00000000",
   247 => x"00000000",
   248 => x"717105ff",
   249 => x"05715351",
   250 => x"020d0400",
   251 => x"00000000",
   252 => x"00000000",
   253 => x"00000000",
   254 => x"00000000",
   255 => x"00000000",
   256 => x"10101010",
   257 => x"10101010",
   258 => x"10101010",
   259 => x"10101010",
   260 => x"10101010",
   261 => x"10101010",
   262 => x"10101010",
   263 => x"10101053",
   264 => x"51047381",
   265 => x"ff067383",
   266 => x"06098105",
   267 => x"83051010",
   268 => x"102b0772",
   269 => x"fc060c51",
   270 => x"51047272",
   271 => x"80728106",
   272 => x"ff050972",
   273 => x"06057110",
   274 => x"52720a10",
   275 => x"0a5372ed",
   276 => x"38515153",
   277 => x"51040000",
   278 => x"800488da",
   279 => x"0488da0b",
   280 => x"8dee0402",
   281 => x"c0050d02",
   282 => x"80c4050b",
   283 => x"0b0ba5a4",
   284 => x"5c5c807c",
   285 => x"7084055e",
   286 => x"08715f5f",
   287 => x"587d7084",
   288 => x"055f0857",
   289 => x"805a7698",
   290 => x"2a77882b",
   291 => x"58557480",
   292 => x"2e81f738",
   293 => x"7c802eb9",
   294 => x"38805d74",
   295 => x"80e42e81",
   296 => x"9f387480",
   297 => x"e42680dc",
   298 => x"387480e3",
   299 => x"2eba38a5",
   300 => x"51989c2d",
   301 => x"7451989c",
   302 => x"2d821858",
   303 => x"811a5a83",
   304 => x"7a25c338",
   305 => x"74ffb638",
   306 => x"7e880c02",
   307 => x"80c0050d",
   308 => x"0474a52e",
   309 => x"09810698",
   310 => x"38810b81",
   311 => x"1b5b5d83",
   312 => x"7a25ffa2",
   313 => x"3889c404",
   314 => x"7b841d71",
   315 => x"08575d54",
   316 => x"7451989c",
   317 => x"2d811881",
   318 => x"1b5b5883",
   319 => x"7a25ff86",
   320 => x"3889c404",
   321 => x"7480f32e",
   322 => x"098106ff",
   323 => x"a2387b84",
   324 => x"1d710870",
   325 => x"545d5d53",
   326 => x"98bd2d80",
   327 => x"0bff1154",
   328 => x"52807225",
   329 => x"ff96387a",
   330 => x"7081055c",
   331 => x"84e02d70",
   332 => x"5255989c",
   333 => x"2d811873",
   334 => x"ff155553",
   335 => x"588aa104",
   336 => x"7b841d71",
   337 => x"087f5c55",
   338 => x"5d528756",
   339 => x"729c2a73",
   340 => x"842b5452",
   341 => x"71802e83",
   342 => x"388159b7",
   343 => x"12547189",
   344 => x"248438b0",
   345 => x"12547892",
   346 => x"38ff1656",
   347 => x"758025dc",
   348 => x"38800bff",
   349 => x"1154528a",
   350 => x"a1047351",
   351 => x"989c2dff",
   352 => x"16567580",
   353 => x"25c6388a",
   354 => x"f1047788",
   355 => x"0c0280c0",
   356 => x"050d04c8",
   357 => x"08880c04",
   358 => x"02fc050d",
   359 => x"80c10b80",
   360 => x"f4f00b85",
   361 => x"802d800b",
   362 => x"80f7880c",
   363 => x"70880c02",
   364 => x"84050d04",
   365 => x"02f8050d",
   366 => x"800b80f4",
   367 => x"f00b84e0",
   368 => x"2d525270",
   369 => x"80c12e9d",
   370 => x"387180f7",
   371 => x"88080780",
   372 => x"f7880c80",
   373 => x"c20b80f4",
   374 => x"f40b8580",
   375 => x"2d70880c",
   376 => x"0288050d",
   377 => x"04810b80",
   378 => x"f7880807",
   379 => x"80f7880c",
   380 => x"80c20b80",
   381 => x"f4f40b85",
   382 => x"802d7088",
   383 => x"0c028805",
   384 => x"0d0402f0",
   385 => x"050d7570",
   386 => x"088a0553",
   387 => x"5380f4f0",
   388 => x"0b84e02d",
   389 => x"517080c1",
   390 => x"2e8c3873",
   391 => x"f0387088",
   392 => x"0c029005",
   393 => x"0d04ff12",
   394 => x"7080f4ec",
   395 => x"0831740c",
   396 => x"880c0290",
   397 => x"050d0402",
   398 => x"ec050d80",
   399 => x"f5980855",
   400 => x"74802e8c",
   401 => x"38767508",
   402 => x"710c80f5",
   403 => x"98085654",
   404 => x"8c155380",
   405 => x"f4ec0852",
   406 => x"8a5195f2",
   407 => x"2d73880c",
   408 => x"0294050d",
   409 => x"0402e805",
   410 => x"0d777008",
   411 => x"5656b053",
   412 => x"80f59808",
   413 => x"5274519d",
   414 => x"e02d850b",
   415 => x"8c170c85",
   416 => x"0b8c160c",
   417 => x"7508750c",
   418 => x"80f59808",
   419 => x"5473802e",
   420 => x"8a387308",
   421 => x"750c80f5",
   422 => x"9808548c",
   423 => x"145380f4",
   424 => x"ec08528a",
   425 => x"5195f22d",
   426 => x"841508ae",
   427 => x"38860b8c",
   428 => x"160c8815",
   429 => x"52881608",
   430 => x"51958c2d",
   431 => x"80f59808",
   432 => x"7008760c",
   433 => x"548c1570",
   434 => x"54548a52",
   435 => x"73085195",
   436 => x"f22d7388",
   437 => x"0c029805",
   438 => x"0d047508",
   439 => x"54b05373",
   440 => x"5275519d",
   441 => x"e02d7388",
   442 => x"0c029805",
   443 => x"0d0402c8",
   444 => x"050d80f4",
   445 => x"840b80f4",
   446 => x"b80c80f4",
   447 => x"bc0b80f5",
   448 => x"980c80f4",
   449 => x"840b80f4",
   450 => x"bc0c800b",
   451 => x"80f4bc0b",
   452 => x"84050c82",
   453 => x"0b80f4bc",
   454 => x"0b88050c",
   455 => x"a80b80f4",
   456 => x"bc0b8c05",
   457 => x"0c9f530b",
   458 => x"0b0ba0a0",
   459 => x"5280f4cc",
   460 => x"519de02d",
   461 => x"9f530b0b",
   462 => x"0ba0c052",
   463 => x"80f6e851",
   464 => x"9de02d8a",
   465 => x"0bb2d00c",
   466 => x"0b0b0ba3",
   467 => x"a05188e3",
   468 => x"2d0b0b0b",
   469 => x"a0e05188",
   470 => x"e32d0b0b",
   471 => x"0ba3a051",
   472 => x"88e32da4",
   473 => x"d008802e",
   474 => x"8499380b",
   475 => x"0b0ba190",
   476 => x"5188e32d",
   477 => x"0b0b0ba3",
   478 => x"a05188e3",
   479 => x"2da4cc08",
   480 => x"520b0b0b",
   481 => x"a1bc5188",
   482 => x"e32dc808",
   483 => x"70a5f00c",
   484 => x"56815880",
   485 => x"0ba4cc08",
   486 => x"2582d838",
   487 => x"02ac055b",
   488 => x"80c10b80",
   489 => x"f4f00b85",
   490 => x"802d810b",
   491 => x"80f7880c",
   492 => x"80c20b80",
   493 => x"f4f40b85",
   494 => x"802d825c",
   495 => x"835a9f53",
   496 => x"0b0b0ba1",
   497 => x"ec5280f4",
   498 => x"f8519de0",
   499 => x"2d815d80",
   500 => x"0b80f4f8",
   501 => x"5380f6e8",
   502 => x"525597a4",
   503 => x"2d880875",
   504 => x"2e098106",
   505 => x"83388155",
   506 => x"7480f788",
   507 => x"0c7b7057",
   508 => x"55748325",
   509 => x"a1387410",
   510 => x"1015fd05",
   511 => x"5e02b805",
   512 => x"fc055383",
   513 => x"52755195",
   514 => x"f22d811c",
   515 => x"705d7057",
   516 => x"55837524",
   517 => x"e1387d54",
   518 => x"7453a5f4",
   519 => x"5280f5a0",
   520 => x"5196842d",
   521 => x"80f59808",
   522 => x"70085757",
   523 => x"b0537652",
   524 => x"75519de0",
   525 => x"2d850b8c",
   526 => x"180c850b",
   527 => x"8c170c76",
   528 => x"08760c80",
   529 => x"f5980855",
   530 => x"74802e8a",
   531 => x"38740876",
   532 => x"0c80f598",
   533 => x"08558c15",
   534 => x"5380f4ec",
   535 => x"08528a51",
   536 => x"95f22d84",
   537 => x"160883e3",
   538 => x"38860b8c",
   539 => x"170c8816",
   540 => x"52881708",
   541 => x"51958c2d",
   542 => x"80f59808",
   543 => x"7008770c",
   544 => x"578c1670",
   545 => x"54558a52",
   546 => x"74085195",
   547 => x"f22d80c1",
   548 => x"0b80f4f4",
   549 => x"0b84e02d",
   550 => x"56567575",
   551 => x"26a53880",
   552 => x"c3527551",
   553 => x"96f02d88",
   554 => x"087d2e82",
   555 => x"ea388116",
   556 => x"7081ff06",
   557 => x"80f4f40b",
   558 => x"84e02d52",
   559 => x"57557476",
   560 => x"27dd387d",
   561 => x"7a7d2935",
   562 => x"705d8a05",
   563 => x"80f4f00b",
   564 => x"84e02d80",
   565 => x"f4ec0859",
   566 => x"57557580",
   567 => x"c12e8386",
   568 => x"3878f738",
   569 => x"811858a4",
   570 => x"cc087825",
   571 => x"fdb238a5",
   572 => x"f00856c8",
   573 => x"087080f4",
   574 => x"b40c7077",
   575 => x"3170a5ec",
   576 => x"0c530b0b",
   577 => x"0ba28c52",
   578 => x"5b88e32d",
   579 => x"a5ec0856",
   580 => x"80f77625",
   581 => x"80f638a4",
   582 => x"cc087077",
   583 => x"87e82935",
   584 => x"a5e40c76",
   585 => x"7187e829",
   586 => x"35a5e80c",
   587 => x"767184b9",
   588 => x"293580f5",
   589 => x"9c0c5a0b",
   590 => x"0b0ba29c",
   591 => x"5188e32d",
   592 => x"a5e40852",
   593 => x"0b0b0ba2",
   594 => x"cc5188e3",
   595 => x"2d0b0b0b",
   596 => x"a2d45188",
   597 => x"e32da5e8",
   598 => x"08520b0b",
   599 => x"0ba2cc51",
   600 => x"88e32d80",
   601 => x"f59c0852",
   602 => x"0b0b0ba3",
   603 => x"845188e3",
   604 => x"2d0b0b0b",
   605 => x"a3a05188",
   606 => x"e32d800b",
   607 => x"880c02b8",
   608 => x"050d040b",
   609 => x"0b0ba3a4",
   610 => x"518ef104",
   611 => x"0b0b0ba3",
   612 => x"d45188e3",
   613 => x"2d0b0b0b",
   614 => x"a48c5188",
   615 => x"e32d0b0b",
   616 => x"0ba3a051",
   617 => x"88e32da5",
   618 => x"ec08a4cc",
   619 => x"08707287",
   620 => x"e82935a5",
   621 => x"e40c7171",
   622 => x"87e82935",
   623 => x"a5e80c71",
   624 => x"7184b929",
   625 => x"3580f59c",
   626 => x"0c5b560b",
   627 => x"0b0ba29c",
   628 => x"5188e32d",
   629 => x"a5e40852",
   630 => x"0b0b0ba2",
   631 => x"cc5188e3",
   632 => x"2d0b0b0b",
   633 => x"a2d45188",
   634 => x"e32da5e8",
   635 => x"08520b0b",
   636 => x"0ba2cc51",
   637 => x"88e32d80",
   638 => x"f59c0852",
   639 => x"0b0b0ba3",
   640 => x"845188e3",
   641 => x"2d0b0b0b",
   642 => x"a3a05188",
   643 => x"e32d800b",
   644 => x"880c02b8",
   645 => x"050d0402",
   646 => x"b805f805",
   647 => x"52805195",
   648 => x"8c2d9f53",
   649 => x"0b0b0ba4",
   650 => x"ac5280f4",
   651 => x"f8519de0",
   652 => x"2d777880",
   653 => x"f4ec0c81",
   654 => x"177081ff",
   655 => x"0680f4f4",
   656 => x"0b84e02d",
   657 => x"5258565a",
   658 => x"91be0476",
   659 => x"0856b053",
   660 => x"75527651",
   661 => x"9de02d80",
   662 => x"c10b80f4",
   663 => x"f40b84e0",
   664 => x"2d565691",
   665 => x"9a04ff15",
   666 => x"7078317c",
   667 => x"0c598059",
   668 => x"91e40402",
   669 => x"f8050d73",
   670 => x"82327009",
   671 => x"81057072",
   672 => x"07802588",
   673 => x"0c525202",
   674 => x"88050d04",
   675 => x"02f4050d",
   676 => x"74767153",
   677 => x"54527182",
   678 => x"2e833883",
   679 => x"5171812e",
   680 => x"9b388172",
   681 => x"26a03871",
   682 => x"822ebc38",
   683 => x"71842eac",
   684 => x"3870730c",
   685 => x"70880c02",
   686 => x"8c050d04",
   687 => x"80e40b80",
   688 => x"f4ec0825",
   689 => x"8c388073",
   690 => x"0c70880c",
   691 => x"028c050d",
   692 => x"0483730c",
   693 => x"70880c02",
   694 => x"8c050d04",
   695 => x"82730c70",
   696 => x"880c028c",
   697 => x"050d0481",
   698 => x"730c7088",
   699 => x"0c028c05",
   700 => x"0d0402fc",
   701 => x"050d7474",
   702 => x"14820571",
   703 => x"0c880c02",
   704 => x"84050d04",
   705 => x"02d8050d",
   706 => x"7b7d7f61",
   707 => x"85127082",
   708 => x"2b751170",
   709 => x"74717084",
   710 => x"05530c5a",
   711 => x"5a5d5b76",
   712 => x"0c7980f8",
   713 => x"180c7986",
   714 => x"12525758",
   715 => x"5a5a7676",
   716 => x"24993876",
   717 => x"b329822b",
   718 => x"79115153",
   719 => x"76737084",
   720 => x"05550c81",
   721 => x"14547574",
   722 => x"25f23876",
   723 => x"81cc2919",
   724 => x"fc110881",
   725 => x"05fc120c",
   726 => x"7a197008",
   727 => x"9fa0130c",
   728 => x"5856850b",
   729 => x"80f4ec0c",
   730 => x"75880c02",
   731 => x"a8050d04",
   732 => x"02f4050d",
   733 => x"02930584",
   734 => x"e02d5180",
   735 => x"02840597",
   736 => x"0584e02d",
   737 => x"54527073",
   738 => x"2e893871",
   739 => x"880c028c",
   740 => x"050d0470",
   741 => x"80f4f00b",
   742 => x"85802d81",
   743 => x"0b880c02",
   744 => x"8c050d04",
   745 => x"02dc050d",
   746 => x"7a7c5956",
   747 => x"820b8319",
   748 => x"55557416",
   749 => x"7084e02d",
   750 => x"7584e02d",
   751 => x"5b515372",
   752 => x"792e80c7",
   753 => x"3880c10b",
   754 => x"81168116",
   755 => x"56565782",
   756 => x"7525df38",
   757 => x"ffa91770",
   758 => x"81ff0655",
   759 => x"59738226",
   760 => x"83388755",
   761 => x"81537680",
   762 => x"d22e9838",
   763 => x"77527551",
   764 => x"9ef92d80",
   765 => x"53728808",
   766 => x"25893887",
   767 => x"1580f4ec",
   768 => x"0c815372",
   769 => x"880c02a4",
   770 => x"050d0472",
   771 => x"80f4f00b",
   772 => x"85802d82",
   773 => x"7525ff9a",
   774 => x"3897d404",
   775 => x"02f8050d",
   776 => x"7352c008",
   777 => x"70882a70",
   778 => x"81065151",
   779 => x"5170802e",
   780 => x"f13871c0",
   781 => x"0c71880c",
   782 => x"0288050d",
   783 => x"0402e805",
   784 => x"0d775675",
   785 => x"70840557",
   786 => x"08538054",
   787 => x"72982a73",
   788 => x"882b5452",
   789 => x"71802ea2",
   790 => x"38c00870",
   791 => x"882a7081",
   792 => x"06515151",
   793 => x"70802ef1",
   794 => x"3871c00c",
   795 => x"81158115",
   796 => x"55558374",
   797 => x"25d63871",
   798 => x"ca387488",
   799 => x"0c029805",
   800 => x"0d049408",
   801 => x"02940cf9",
   802 => x"3d0d800b",
   803 => x"9408fc05",
   804 => x"0c940888",
   805 => x"05088025",
   806 => x"ab389408",
   807 => x"88050830",
   808 => x"94088805",
   809 => x"0c800b94",
   810 => x"08f4050c",
   811 => x"9408fc05",
   812 => x"08883881",
   813 => x"0b9408f4",
   814 => x"050c9408",
   815 => x"f4050894",
   816 => x"08fc050c",
   817 => x"94088c05",
   818 => x"088025ab",
   819 => x"3894088c",
   820 => x"05083094",
   821 => x"088c050c",
   822 => x"800b9408",
   823 => x"f0050c94",
   824 => x"08fc0508",
   825 => x"8838810b",
   826 => x"9408f005",
   827 => x"0c9408f0",
   828 => x"05089408",
   829 => x"fc050c80",
   830 => x"5394088c",
   831 => x"05085294",
   832 => x"08880508",
   833 => x"5181a73f",
   834 => x"88087094",
   835 => x"08f8050c",
   836 => x"549408fc",
   837 => x"0508802e",
   838 => x"8c389408",
   839 => x"f8050830",
   840 => x"9408f805",
   841 => x"0c9408f8",
   842 => x"05087088",
   843 => x"0c54893d",
   844 => x"0d940c04",
   845 => x"94080294",
   846 => x"0cfb3d0d",
   847 => x"800b9408",
   848 => x"fc050c94",
   849 => x"08880508",
   850 => x"80259338",
   851 => x"94088805",
   852 => x"08309408",
   853 => x"88050c81",
   854 => x"0b9408fc",
   855 => x"050c9408",
   856 => x"8c050880",
   857 => x"258c3894",
   858 => x"088c0508",
   859 => x"3094088c",
   860 => x"050c8153",
   861 => x"94088c05",
   862 => x"08529408",
   863 => x"88050851",
   864 => x"ad3f8808",
   865 => x"709408f8",
   866 => x"050c5494",
   867 => x"08fc0508",
   868 => x"802e8c38",
   869 => x"9408f805",
   870 => x"08309408",
   871 => x"f8050c94",
   872 => x"08f80508",
   873 => x"70880c54",
   874 => x"873d0d94",
   875 => x"0c049408",
   876 => x"02940cfd",
   877 => x"3d0d810b",
   878 => x"9408fc05",
   879 => x"0c800b94",
   880 => x"08f8050c",
   881 => x"94088c05",
   882 => x"08940888",
   883 => x"050827ac",
   884 => x"389408fc",
   885 => x"0508802e",
   886 => x"a338800b",
   887 => x"94088c05",
   888 => x"08249938",
   889 => x"94088c05",
   890 => x"08109408",
   891 => x"8c050c94",
   892 => x"08fc0508",
   893 => x"109408fc",
   894 => x"050cc939",
   895 => x"9408fc05",
   896 => x"08802e80",
   897 => x"c9389408",
   898 => x"8c050894",
   899 => x"08880508",
   900 => x"26a13894",
   901 => x"08880508",
   902 => x"94088c05",
   903 => x"08319408",
   904 => x"88050c94",
   905 => x"08f80508",
   906 => x"9408fc05",
   907 => x"08079408",
   908 => x"f8050c94",
   909 => x"08fc0508",
   910 => x"812a9408",
   911 => x"fc050c94",
   912 => x"088c0508",
   913 => x"812a9408",
   914 => x"8c050cff",
   915 => x"af399408",
   916 => x"90050880",
   917 => x"2e8f3894",
   918 => x"08880508",
   919 => x"709408f4",
   920 => x"050c518d",
   921 => x"399408f8",
   922 => x"05087094",
   923 => x"08f4050c",
   924 => x"519408f4",
   925 => x"0508880c",
   926 => x"853d0d94",
   927 => x"0c049408",
   928 => x"02940cff",
   929 => x"3d0d800b",
   930 => x"9408fc05",
   931 => x"0c940888",
   932 => x"05088106",
   933 => x"ff117009",
   934 => x"7094088c",
   935 => x"05080694",
   936 => x"08fc0508",
   937 => x"119408fc",
   938 => x"050c9408",
   939 => x"88050881",
   940 => x"2a940888",
   941 => x"050c9408",
   942 => x"8c050810",
   943 => x"94088c05",
   944 => x"0c515151",
   945 => x"51940888",
   946 => x"0508802e",
   947 => x"8438ffbd",
   948 => x"399408fc",
   949 => x"05087088",
   950 => x"0c51833d",
   951 => x"0d940c04",
   952 => x"fc3d0d76",
   953 => x"70797b55",
   954 => x"5555558f",
   955 => x"72278c38",
   956 => x"72750783",
   957 => x"06517080",
   958 => x"2ea738ff",
   959 => x"125271ff",
   960 => x"2e983872",
   961 => x"70810554",
   962 => x"33747081",
   963 => x"055634ff",
   964 => x"125271ff",
   965 => x"2e098106",
   966 => x"ea387488",
   967 => x"0c863d0d",
   968 => x"04745172",
   969 => x"70840554",
   970 => x"08717084",
   971 => x"05530c72",
   972 => x"70840554",
   973 => x"08717084",
   974 => x"05530c72",
   975 => x"70840554",
   976 => x"08717084",
   977 => x"05530c72",
   978 => x"70840554",
   979 => x"08717084",
   980 => x"05530cf0",
   981 => x"1252718f",
   982 => x"26c93883",
   983 => x"72279538",
   984 => x"72708405",
   985 => x"54087170",
   986 => x"8405530c",
   987 => x"fc125271",
   988 => x"8326ed38",
   989 => x"7054ff83",
   990 => x"39fb3d0d",
   991 => x"77797072",
   992 => x"07830653",
   993 => x"54527093",
   994 => x"38717373",
   995 => x"08545654",
   996 => x"7173082e",
   997 => x"80c43873",
   998 => x"75545271",
   999 => x"337081ff",
  1000 => x"06525470",
  1001 => x"802e9d38",
  1002 => x"72335570",
  1003 => x"752e0981",
  1004 => x"06953881",
  1005 => x"12811471",
  1006 => x"337081ff",
  1007 => x"06545654",
  1008 => x"5270e538",
  1009 => x"72335573",
  1010 => x"81ff0675",
  1011 => x"81ff0671",
  1012 => x"7131880c",
  1013 => x"5252873d",
  1014 => x"0d047109",
  1015 => x"70f7fbfd",
  1016 => x"ff140670",
  1017 => x"f8848281",
  1018 => x"80065151",
  1019 => x"51709738",
  1020 => x"84148416",
  1021 => x"71085456",
  1022 => x"54717508",
  1023 => x"2edc3873",
  1024 => x"755452ff",
  1025 => x"9639800b",
  1026 => x"880c873d",
  1027 => x"0d040000",
  1028 => x"00ffffff",
  1029 => x"ff00ffff",
  1030 => x"ffff00ff",
  1031 => x"ffffff00",
  1032 => x"44485259",
  1033 => x"53544f4e",
  1034 => x"45205052",
  1035 => x"4f475241",
  1036 => x"4d2c2053",
  1037 => x"4f4d4520",
  1038 => x"53545249",
  1039 => x"4e470000",
  1040 => x"44485259",
  1041 => x"53544f4e",
  1042 => x"45205052",
  1043 => x"4f475241",
  1044 => x"4d2c2031",
  1045 => x"27535420",
  1046 => x"53545249",
  1047 => x"4e470000",
  1048 => x"44687279",
  1049 => x"73746f6e",
  1050 => x"65204265",
  1051 => x"6e63686d",
  1052 => x"61726b2c",
  1053 => x"20566572",
  1054 => x"73696f6e",
  1055 => x"20322e31",
  1056 => x"20284c61",
  1057 => x"6e677561",
  1058 => x"67653a20",
  1059 => x"43290a00",
  1060 => x"50726f67",
  1061 => x"72616d20",
  1062 => x"636f6d70",
  1063 => x"696c6564",
  1064 => x"20776974",
  1065 => x"68202772",
  1066 => x"65676973",
  1067 => x"74657227",
  1068 => x"20617474",
  1069 => x"72696275",
  1070 => x"74650a00",
  1071 => x"45786563",
  1072 => x"7574696f",
  1073 => x"6e207374",
  1074 => x"61727473",
  1075 => x"2c202564",
  1076 => x"2072756e",
  1077 => x"73207468",
  1078 => x"726f7567",
  1079 => x"68204468",
  1080 => x"72797374",
  1081 => x"6f6e650a",
  1082 => x"00000000",
  1083 => x"44485259",
  1084 => x"53544f4e",
  1085 => x"45205052",
  1086 => x"4f475241",
  1087 => x"4d2c2032",
  1088 => x"274e4420",
  1089 => x"53545249",
  1090 => x"4e470000",
  1091 => x"55736572",
  1092 => x"2074696d",
  1093 => x"653a2025",
  1094 => x"640a0000",
  1095 => x"4d696372",
  1096 => x"6f736563",
  1097 => x"6f6e6473",
  1098 => x"20666f72",
  1099 => x"206f6e65",
  1100 => x"2072756e",
  1101 => x"20746872",
  1102 => x"6f756768",
  1103 => x"20446872",
  1104 => x"7973746f",
  1105 => x"6e653a20",
  1106 => x"00000000",
  1107 => x"2564200a",
  1108 => x"00000000",
  1109 => x"44687279",
  1110 => x"73746f6e",
  1111 => x"65732070",
  1112 => x"65722053",
  1113 => x"65636f6e",
  1114 => x"643a2020",
  1115 => x"20202020",
  1116 => x"20202020",
  1117 => x"20202020",
  1118 => x"20202020",
  1119 => x"20202020",
  1120 => x"00000000",
  1121 => x"56415820",
  1122 => x"4d495053",
  1123 => x"20726174",
  1124 => x"696e6720",
  1125 => x"2a203130",
  1126 => x"3030203d",
  1127 => x"20256420",
  1128 => x"0a000000",
  1129 => x"50726f67",
  1130 => x"72616d20",
  1131 => x"636f6d70",
  1132 => x"696c6564",
  1133 => x"20776974",
  1134 => x"686f7574",
  1135 => x"20277265",
  1136 => x"67697374",
  1137 => x"65722720",
  1138 => x"61747472",
  1139 => x"69627574",
  1140 => x"650a0000",
  1141 => x"4d656173",
  1142 => x"75726564",
  1143 => x"2074696d",
  1144 => x"6520746f",
  1145 => x"6f20736d",
  1146 => x"616c6c20",
  1147 => x"746f206f",
  1148 => x"62746169",
  1149 => x"6e206d65",
  1150 => x"616e696e",
  1151 => x"6766756c",
  1152 => x"20726573",
  1153 => x"756c7473",
  1154 => x"0a000000",
  1155 => x"506c6561",
  1156 => x"73652069",
  1157 => x"6e637265",
  1158 => x"61736520",
  1159 => x"6e756d62",
  1160 => x"6572206f",
  1161 => x"66207275",
  1162 => x"6e730a00",
  1163 => x"44485259",
  1164 => x"53544f4e",
  1165 => x"45205052",
  1166 => x"4f475241",
  1167 => x"4d2c2033",
  1168 => x"27524420",
  1169 => x"53545249",
  1170 => x"4e470000",
  1171 => x"000061a8",
  1172 => x"00000000",
	others => x"00000000"
);

begin

process (clk)
begin
	if (clk'event and clk = '1') then
		if (from_zpu.memAWriteEnable = '1') and (from_zpu.memBWriteEnable = '1') and (from_zpu.memAAddr=from_zpu.memBAddr) and (from_zpu.memAWrite/=from_zpu.memBWrite) then
			report "write collision" severity failure;
		end if;
	
		if (from_zpu.memAWriteEnable = '1') then
			ram(to_integer(unsigned(from_zpu.memAAddr(maxAddrBit downto 2)))) := from_zpu.memAWrite;
			to_zpu.memARead <= from_zpu.memAWrite;
		else
			to_zpu.memARead <= ram(to_integer(unsigned(from_zpu.memAAddr(maxAddrBit downto 2))));
		end if;
	end if;
end process;

process (clk)
begin
	if (clk'event and clk = '1') then
		if (from_zpu.memBWriteEnable = '1') then
			ram(to_integer(unsigned(from_zpu.memBAddr(maxAddrBit downto 2)))) := from_zpu.memBWrite;
			to_zpu.memBRead <= from_zpu.memBWrite;
		else
			to_zpu.memBRead <= ram(to_integer(unsigned(from_zpu.memBAddr(maxAddrBit downto 2))));
		end if;
	end if;
end process;


end arch;

