-- ZPU
--
-- Copyright 2004-2008 oharboe - �yvind Harboe - oyvind.harboe@zylin.com
-- Modified by Alastair M. Robinson for the ZPUFlex project.
--
-- The FreeBSD license
-- 
-- Redistribution and use in source and binary forms, with or without
-- modification, are permitted provided that the following conditions
-- are met:
-- 
-- 1. Redistributions of source code must retain the above copyright
--    notice, this list of conditions and the following disclaimer.
-- 2. Redistributions in binary form must reproduce the above
--    copyright notice, this list of conditions and the following
--    disclaimer in the documentation and/or other materials
--    provided with the distribution.
-- 
-- THIS SOFTWARE IS PROVIDED BY THE ZPU PROJECT ``AS IS'' AND ANY
-- EXPRESS OR IMPLIED WARRANTIES, INCLUDING, BUT NOT LIMITED TO,
-- THE IMPLIED WARRANTIES OF MERCHANTABILITY AND FITNESS FOR A
-- PARTICULAR PURPOSE ARE DISCLAIMED. IN NO EVENT SHALL THE
-- ZPU PROJECT OR CONTRIBUTORS BE LIABLE FOR ANY DIRECT,
-- INDIRECT, INCIDENTAL, SPECIAL, EXEMPLARY, OR CONSEQUENTIAL DAMAGES
-- (INCLUDING, BUT NOT LIMITED TO, PROCUREMENT OF SUBSTITUTE GOODS
-- OR SERVICES; LOSS OF USE, DATA, OR PROFITS; OR BUSINESS INTERRUPTION)
-- HOWEVER CAUSED AND ON ANY THEORY OF LIABILITY, WHETHER IN CONTRACT,
-- STRICT LIABILITY, OR TORT (INCLUDING NEGLIGENCE OR OTHERWISE)
-- ARISING IN ANY WAY OUT OF THE USE OF THIS SOFTWARE, EVEN IF
-- ADVISED OF THE POSSIBILITY OF SUCH DAMAGE.
-- 
-- The views and conclusions contained in the software and documentation
-- are those of the authors and should not be interpreted as representing
-- official policies, either expressed or implied, of the ZPU Project.

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;


library work;
use work.zpupkg.all;

entity SDBootstrap_ROM is
generic
	(
		maxAddrBitBRAM : integer := maxAddrBitBRAMLimit -- Specify your actual ROM size to save LEs and unnecessary block RAM usage.
	);
port (
	clk : in std_logic;
	areset : in std_logic := '0';
	from_zpu : in ZPU_ToROM;
	to_zpu : out ZPU_FromROM
);
end SDBootstrap_ROM;

architecture arch of SDBootstrap_ROM is

type ram_type is array(natural range 0 to ((2**(maxAddrBitBRAM+1))/4)-1) of std_logic_vector(wordSize-1 downto 0);

shared variable ram : ram_type :=
(
     0 => x"84808080",
     1 => x"ee040000",
     2 => x"00000000",
     3 => x"84808080",
     4 => x"88080d80",
     5 => x"04848080",
     6 => x"80950471",
     7 => x"fd060872",
     8 => x"83060981",
     9 => x"05820583",
    10 => x"2b2a83ff",
    11 => x"ff065204",
    12 => x"71fc0608",
    13 => x"72830609",
    14 => x"81058305",
    15 => x"1010102a",
    16 => x"81ff0652",
    17 => x"0471fc06",
    18 => x"08848080",
    19 => x"a1c87383",
    20 => x"06101005",
    21 => x"08067381",
    22 => x"ff067383",
    23 => x"06098105",
    24 => x"83051010",
    25 => x"102b0772",
    26 => x"fc060c51",
    27 => x"51040284",
    28 => x"05848080",
    29 => x"80880c84",
    30 => x"80808095",
    31 => x"0b848080",
    32 => x"8ed10400",
    33 => x"02ec050d",
    34 => x"76538055",
    35 => x"7275258e",
    36 => x"38ad5184",
    37 => x"808084b2",
    38 => x"2d720981",
    39 => x"05537280",
    40 => x"2ebe3887",
    41 => x"54729c2a",
    42 => x"73842b54",
    43 => x"5271802e",
    44 => x"83388155",
    45 => x"8972258a",
    46 => x"38b71252",
    47 => x"84808081",
    48 => x"c504b012",
    49 => x"5274802e",
    50 => x"89387151",
    51 => x"84808084",
    52 => x"b22dff14",
    53 => x"54738025",
    54 => x"cc388480",
    55 => x"8081e804",
    56 => x"b0518480",
    57 => x"8084b22d",
    58 => x"800b83ff",
    59 => x"e0800c02",
    60 => x"94050d04",
    61 => x"02c0050d",
    62 => x"0280c405",
    63 => x"57807078",
    64 => x"7084055a",
    65 => x"0872415f",
    66 => x"5d587c70",
    67 => x"84055e08",
    68 => x"5a805b79",
    69 => x"982a7a88",
    70 => x"2b5b5675",
    71 => x"8938775f",
    72 => x"84808084",
    73 => x"a6047d80",
    74 => x"2e81d338",
    75 => x"805e7580",
    76 => x"e42e8a38",
    77 => x"7580f82e",
    78 => x"09810689",
    79 => x"38768418",
    80 => x"71085e58",
    81 => x"547580e4",
    82 => x"2ea63875",
    83 => x"80e4268e",
    84 => x"387580e3",
    85 => x"2e80d938",
    86 => x"84808083",
    87 => x"be047580",
    88 => x"f32eb538",
    89 => x"7580f82e",
    90 => x"8f388480",
    91 => x"8083be04",
    92 => x"8a538480",
    93 => x"8082fa04",
    94 => x"905383ff",
    95 => x"e0e0527b",
    96 => x"51848080",
    97 => x"81842d83",
    98 => x"ffe08008",
    99 => x"83ffe0e0",
   100 => x"5a558480",
   101 => x"8083d704",
   102 => x"76841871",
   103 => x"0870545b",
   104 => x"58548480",
   105 => x"8084d62d",
   106 => x"80558480",
   107 => x"8083d704",
   108 => x"76841871",
   109 => x"08585854",
   110 => x"84808084",
   111 => x"8e04a551",
   112 => x"84808084",
   113 => x"b22d7551",
   114 => x"84808084",
   115 => x"b22d8218",
   116 => x"58848080",
   117 => x"84990474",
   118 => x"ff165654",
   119 => x"807425b9",
   120 => x"38787081",
   121 => x"055a8480",
   122 => x"8080b02d",
   123 => x"70525684",
   124 => x"808084b2",
   125 => x"2d811858",
   126 => x"84808083",
   127 => x"d70475a5",
   128 => x"2e098106",
   129 => x"8938815e",
   130 => x"84808084",
   131 => x"99047551",
   132 => x"84808084",
   133 => x"b22d8118",
   134 => x"58811b5b",
   135 => x"837b25fd",
   136 => x"f23875fd",
   137 => x"e5387e83",
   138 => x"ffe0800c",
   139 => x"0280c005",
   140 => x"0d0402f8",
   141 => x"050d7352",
   142 => x"c0087088",
   143 => x"2a708106",
   144 => x"51515170",
   145 => x"802ef138",
   146 => x"71c00c71",
   147 => x"83ffe080",
   148 => x"0c028805",
   149 => x"0d0402e8",
   150 => x"050d8078",
   151 => x"57557570",
   152 => x"84055708",
   153 => x"53805472",
   154 => x"982a7388",
   155 => x"2b545271",
   156 => x"802ea238",
   157 => x"c0087088",
   158 => x"2a708106",
   159 => x"51515170",
   160 => x"802ef138",
   161 => x"71c00c81",
   162 => x"15811555",
   163 => x"55837425",
   164 => x"d63871ca",
   165 => x"387483ff",
   166 => x"e0800c02",
   167 => x"98050d04",
   168 => x"02f4050d",
   169 => x"d45281ff",
   170 => x"720c7108",
   171 => x"5381ff72",
   172 => x"0c72882b",
   173 => x"83fe8006",
   174 => x"72087081",
   175 => x"ff065152",
   176 => x"5381ff72",
   177 => x"0c727107",
   178 => x"882b7208",
   179 => x"7081ff06",
   180 => x"51525381",
   181 => x"ff720c72",
   182 => x"7107882b",
   183 => x"72087081",
   184 => x"ff067207",
   185 => x"83ffe080",
   186 => x"0c525302",
   187 => x"8c050d04",
   188 => x"02f4050d",
   189 => x"74767181",
   190 => x"ff06d40c",
   191 => x"535383ff",
   192 => x"f1a00885",
   193 => x"3871892b",
   194 => x"5271982a",
   195 => x"d40c7190",
   196 => x"2a7081ff",
   197 => x"06d40c51",
   198 => x"71882a70",
   199 => x"81ff06d4",
   200 => x"0c517181",
   201 => x"ff06d40c",
   202 => x"72902a70",
   203 => x"81ff06d4",
   204 => x"0c51d408",
   205 => x"7081ff06",
   206 => x"515182b8",
   207 => x"bf527081",
   208 => x"ff2e0981",
   209 => x"06943881",
   210 => x"ff0bd40c",
   211 => x"d4087081",
   212 => x"ff06ff14",
   213 => x"54515171",
   214 => x"e5387083",
   215 => x"ffe0800c",
   216 => x"028c050d",
   217 => x"0402fc05",
   218 => x"0d81c751",
   219 => x"81ff0bd4",
   220 => x"0cff1151",
   221 => x"708025f4",
   222 => x"38028405",
   223 => x"0d0402f0",
   224 => x"050d8480",
   225 => x"8086e52d",
   226 => x"819c9f53",
   227 => x"805287fc",
   228 => x"80f75184",
   229 => x"808085f0",
   230 => x"2d83ffe0",
   231 => x"80085483",
   232 => x"ffe08008",
   233 => x"812e0981",
   234 => x"06ae3881",
   235 => x"ff0bd40c",
   236 => x"820a5284",
   237 => x"9c80e951",
   238 => x"84808085",
   239 => x"f02d83ff",
   240 => x"e080088e",
   241 => x"3881ff0b",
   242 => x"d40c7353",
   243 => x"84808087",
   244 => x"df048480",
   245 => x"8086e52d",
   246 => x"ff135372",
   247 => x"ffae3872",
   248 => x"83ffe080",
   249 => x"0c029005",
   250 => x"0d0402f4",
   251 => x"050d81ff",
   252 => x"0bd40c84",
   253 => x"8080a1d8",
   254 => x"51848080",
   255 => x"84d62d93",
   256 => x"53805287",
   257 => x"fc80c151",
   258 => x"84808085",
   259 => x"f02d83ff",
   260 => x"e080088e",
   261 => x"3881ff0b",
   262 => x"d40c8153",
   263 => x"84808088",
   264 => x"ae048480",
   265 => x"8086e52d",
   266 => x"ff135372",
   267 => x"d4387283",
   268 => x"ffe0800c",
   269 => x"028c050d",
   270 => x"0402f005",
   271 => x"0d848080",
   272 => x"86e52d83",
   273 => x"aa52849c",
   274 => x"80c85184",
   275 => x"808085f0",
   276 => x"2d83ffe0",
   277 => x"800883ff",
   278 => x"e0800853",
   279 => x"848080a1",
   280 => x"e4525384",
   281 => x"808081f4",
   282 => x"2d72812e",
   283 => x"098106a9",
   284 => x"38848080",
   285 => x"85a02d83",
   286 => x"ffe08008",
   287 => x"83ffff06",
   288 => x"537283aa",
   289 => x"2ebb3883",
   290 => x"ffe08008",
   291 => x"52848080",
   292 => x"a1fc5184",
   293 => x"808081f4",
   294 => x"2d848080",
   295 => x"87ea2d84",
   296 => x"808089b9",
   297 => x"04815484",
   298 => x"80808ae4",
   299 => x"04848080",
   300 => x"a2945184",
   301 => x"808081f4",
   302 => x"2d805484",
   303 => x"80808ae4",
   304 => x"0481ff0b",
   305 => x"d40cb153",
   306 => x"84808086",
   307 => x"fe2d83ff",
   308 => x"e0800880",
   309 => x"2e80fe38",
   310 => x"805287fc",
   311 => x"80fa5184",
   312 => x"808085f0",
   313 => x"2d83ffe0",
   314 => x"800880d7",
   315 => x"3883ffe0",
   316 => x"80085284",
   317 => x"8080a2b0",
   318 => x"51848080",
   319 => x"81f42d81",
   320 => x"ff0bd40c",
   321 => x"d4087081",
   322 => x"ff067054",
   323 => x"848080a2",
   324 => x"bc535153",
   325 => x"84808081",
   326 => x"f42d81ff",
   327 => x"0bd40c81",
   328 => x"ff0bd40c",
   329 => x"81ff0bd4",
   330 => x"0c81ff0b",
   331 => x"d40c7286",
   332 => x"2a708106",
   333 => x"70565153",
   334 => x"72802ea8",
   335 => x"38848080",
   336 => x"89a50483",
   337 => x"ffe08008",
   338 => x"52848080",
   339 => x"a2b05184",
   340 => x"808081f4",
   341 => x"2d72822e",
   342 => x"fed338ff",
   343 => x"135372fe",
   344 => x"e7387254",
   345 => x"7383ffe0",
   346 => x"800c0290",
   347 => x"050d0402",
   348 => x"f4050d81",
   349 => x"0b83fff1",
   350 => x"a00cd008",
   351 => x"708f2a70",
   352 => x"81065151",
   353 => x"5372f338",
   354 => x"72d00c84",
   355 => x"808086e5",
   356 => x"2d848080",
   357 => x"a2cc5184",
   358 => x"808084d6",
   359 => x"2dd00870",
   360 => x"8f2a7081",
   361 => x"06515153",
   362 => x"72f33881",
   363 => x"0bd00c87",
   364 => x"53805284",
   365 => x"d480c051",
   366 => x"84808085",
   367 => x"f02d83ff",
   368 => x"e0800881",
   369 => x"2e973872",
   370 => x"822e0981",
   371 => x"06893880",
   372 => x"53848080",
   373 => x"8c9704ff",
   374 => x"135372d5",
   375 => x"38848080",
   376 => x"88b92d83",
   377 => x"ffe08008",
   378 => x"83fff1a0",
   379 => x"0c815287",
   380 => x"fc80d051",
   381 => x"84808085",
   382 => x"f02d81ff",
   383 => x"0bd40cd0",
   384 => x"08708f2a",
   385 => x"70810651",
   386 => x"515372f3",
   387 => x"3872d00c",
   388 => x"81ff0bd4",
   389 => x"0c815372",
   390 => x"83ffe080",
   391 => x"0c028c05",
   392 => x"0d04800b",
   393 => x"83ffe080",
   394 => x"0c0402e0",
   395 => x"050d797b",
   396 => x"57578058",
   397 => x"81ff0bd4",
   398 => x"0cd00870",
   399 => x"8f2a7081",
   400 => x"06515154",
   401 => x"73f33882",
   402 => x"810bd00c",
   403 => x"81ff0bd4",
   404 => x"0c765287",
   405 => x"fc80d151",
   406 => x"84808085",
   407 => x"f02d80db",
   408 => x"c6df5583",
   409 => x"ffe08008",
   410 => x"802e9b38",
   411 => x"83ffe080",
   412 => x"08537652",
   413 => x"848080a2",
   414 => x"d8518480",
   415 => x"8081f42d",
   416 => x"8480808d",
   417 => x"dc0481ff",
   418 => x"0bd40cd4",
   419 => x"087081ff",
   420 => x"06515473",
   421 => x"81fe2e09",
   422 => x"8106a538",
   423 => x"80ff5484",
   424 => x"808085a0",
   425 => x"2d83ffe0",
   426 => x"80087670",
   427 => x"8405580c",
   428 => x"ff145473",
   429 => x"8025e838",
   430 => x"81588480",
   431 => x"808dc604",
   432 => x"ff155574",
   433 => x"c13881ff",
   434 => x"0bd40cd0",
   435 => x"08708f2a",
   436 => x"70810651",
   437 => x"515473f3",
   438 => x"3873d00c",
   439 => x"7783ffe0",
   440 => x"800c02a0",
   441 => x"050d0402",
   442 => x"f4050d74",
   443 => x"70882a83",
   444 => x"fe800670",
   445 => x"72982a07",
   446 => x"72882b87",
   447 => x"fc808006",
   448 => x"73982b81",
   449 => x"f00a0671",
   450 => x"73070783",
   451 => x"ffe0800c",
   452 => x"56515351",
   453 => x"028c050d",
   454 => x"0402f805",
   455 => x"0d028e05",
   456 => x"84808080",
   457 => x"b02d7488",
   458 => x"2b077083",
   459 => x"ffff0683",
   460 => x"ffe0800c",
   461 => x"51028805",
   462 => x"0d0402f8",
   463 => x"050d7370",
   464 => x"902b7190",
   465 => x"2a0783ff",
   466 => x"e0800c52",
   467 => x"0288050d",
   468 => x"0402ec05",
   469 => x"0d800bfc",
   470 => x"800c8480",
   471 => x"80a2f851",
   472 => x"84808084",
   473 => x"d62d8480",
   474 => x"808aef2d",
   475 => x"83ffe080",
   476 => x"08802e82",
   477 => x"86388480",
   478 => x"80a39051",
   479 => x"84808084",
   480 => x"d62d8480",
   481 => x"8091df2d",
   482 => x"83ffe1a0",
   483 => x"52848080",
   484 => x"a3a85184",
   485 => x"80809ee0",
   486 => x"2d83ffe0",
   487 => x"8008802e",
   488 => x"81cd3883",
   489 => x"ffe1a00b",
   490 => x"848080a3",
   491 => x"b4525484",
   492 => x"808084d6",
   493 => x"2d805573",
   494 => x"70810555",
   495 => x"84808080",
   496 => x"b02d5372",
   497 => x"a02e80e6",
   498 => x"3872c00c",
   499 => x"72a32e81",
   500 => x"84387280",
   501 => x"c72e0981",
   502 => x"068d3884",
   503 => x"8080808c",
   504 => x"2d848080",
   505 => x"90890472",
   506 => x"8a2e0981",
   507 => x"068d3884",
   508 => x"80808095",
   509 => x"2d848080",
   510 => x"90890472",
   511 => x"80cc2e09",
   512 => x"81068638",
   513 => x"83ffe1a0",
   514 => x"547281df",
   515 => x"06f00570",
   516 => x"81ff0651",
   517 => x"53b87327",
   518 => x"8938ef13",
   519 => x"7081ff06",
   520 => x"51537484",
   521 => x"2b730755",
   522 => x"8480808f",
   523 => x"b70472a3",
   524 => x"2ea33873",
   525 => x"70810555",
   526 => x"84808080",
   527 => x"b02d5372",
   528 => x"a02ef038",
   529 => x"ff147553",
   530 => x"70525484",
   531 => x"80809ee0",
   532 => x"2d74fc80",
   533 => x"0c737081",
   534 => x"05558480",
   535 => x"8080b02d",
   536 => x"53728a2e",
   537 => x"098106ed",
   538 => x"38848080",
   539 => x"8fb50484",
   540 => x"8080a3c8",
   541 => x"51848080",
   542 => x"84d62d84",
   543 => x"8080a3e4",
   544 => x"51848080",
   545 => x"84d62d80",
   546 => x"0b83ffe0",
   547 => x"800c0294",
   548 => x"050d0402",
   549 => x"e8050d77",
   550 => x"797b5855",
   551 => x"55805372",
   552 => x"7625af38",
   553 => x"74708105",
   554 => x"56848080",
   555 => x"80b02d74",
   556 => x"70810556",
   557 => x"84808080",
   558 => x"b02d5252",
   559 => x"71712e89",
   560 => x"38815184",
   561 => x"808091d4",
   562 => x"04811353",
   563 => x"84808091",
   564 => x"9f048051",
   565 => x"7083ffe0",
   566 => x"800c0298",
   567 => x"050d0402",
   568 => x"d8050dff",
   569 => x"0b83fff5",
   570 => x"cc0c800b",
   571 => x"83fff5e0",
   572 => x"0c848080",
   573 => x"a3f05184",
   574 => x"808084d6",
   575 => x"2d83fff1",
   576 => x"b8528051",
   577 => x"8480808c",
   578 => x"aa2d83ff",
   579 => x"e0800854",
   580 => x"83ffe080",
   581 => x"08953884",
   582 => x"8080a480",
   583 => x"51848080",
   584 => x"84d62d73",
   585 => x"55848080",
   586 => x"9a950484",
   587 => x"8080a494",
   588 => x"51848080",
   589 => x"84d62d80",
   590 => x"56810b83",
   591 => x"fff1ac0c",
   592 => x"88538480",
   593 => x"80a4ac52",
   594 => x"83fff1ee",
   595 => x"51848080",
   596 => x"91932d83",
   597 => x"ffe08008",
   598 => x"762e0981",
   599 => x"068b3883",
   600 => x"ffe08008",
   601 => x"83fff1ac",
   602 => x"0c885384",
   603 => x"8080a4b8",
   604 => x"5283fff2",
   605 => x"8a518480",
   606 => x"8091932d",
   607 => x"83ffe080",
   608 => x"088b3883",
   609 => x"ffe08008",
   610 => x"83fff1ac",
   611 => x"0c83fff1",
   612 => x"ac085284",
   613 => x"8080a4c4",
   614 => x"51848080",
   615 => x"81f42d83",
   616 => x"fff1ac08",
   617 => x"802e81cb",
   618 => x"3883fff4",
   619 => x"fe0b8480",
   620 => x"8080b02d",
   621 => x"83fff4ff",
   622 => x"0b848080",
   623 => x"80b02d71",
   624 => x"982b7190",
   625 => x"2b0783ff",
   626 => x"f5800b84",
   627 => x"808080b0",
   628 => x"2d70882b",
   629 => x"720783ff",
   630 => x"f5810b84",
   631 => x"808080b0",
   632 => x"2d710783",
   633 => x"fff5b60b",
   634 => x"84808080",
   635 => x"b02d83ff",
   636 => x"f5b70b84",
   637 => x"808080b0",
   638 => x"2d71882b",
   639 => x"07535f54",
   640 => x"525a5657",
   641 => x"557381ab",
   642 => x"aa2e0981",
   643 => x"06953875",
   644 => x"51848080",
   645 => x"8de72d83",
   646 => x"ffe08008",
   647 => x"56848080",
   648 => x"94bc0473",
   649 => x"82d4d52e",
   650 => x"93388480",
   651 => x"80a4d851",
   652 => x"84808084",
   653 => x"d62d8480",
   654 => x"8096c804",
   655 => x"75528480",
   656 => x"80a4f851",
   657 => x"84808081",
   658 => x"f42d83ff",
   659 => x"f1b85275",
   660 => x"51848080",
   661 => x"8caa2d83",
   662 => x"ffe08008",
   663 => x"5583ffe0",
   664 => x"8008802e",
   665 => x"85af3884",
   666 => x"8080a590",
   667 => x"51848080",
   668 => x"84d62d84",
   669 => x"8080a5b8",
   670 => x"51848080",
   671 => x"81f42d88",
   672 => x"53848080",
   673 => x"a4b85283",
   674 => x"fff28a51",
   675 => x"84808091",
   676 => x"932d83ff",
   677 => x"e080088e",
   678 => x"38810b83",
   679 => x"fff5e00c",
   680 => x"84808095",
   681 => x"d4048853",
   682 => x"848080a4",
   683 => x"ac5283ff",
   684 => x"f1ee5184",
   685 => x"80809193",
   686 => x"2d83ffe0",
   687 => x"8008802e",
   688 => x"93388480",
   689 => x"80a5d051",
   690 => x"84808081",
   691 => x"f42d8480",
   692 => x"8096c804",
   693 => x"83fff5b6",
   694 => x"0b848080",
   695 => x"80b02d54",
   696 => x"7380d52e",
   697 => x"09810680",
   698 => x"df3883ff",
   699 => x"f5b70b84",
   700 => x"808080b0",
   701 => x"2d547381",
   702 => x"aa2e0981",
   703 => x"0680c938",
   704 => x"800b83ff",
   705 => x"f1b80b84",
   706 => x"808080b0",
   707 => x"2d565474",
   708 => x"81e92e83",
   709 => x"38815474",
   710 => x"81eb2e8c",
   711 => x"38805573",
   712 => x"752e0981",
   713 => x"0683ee38",
   714 => x"83fff1c3",
   715 => x"0b848080",
   716 => x"80b02d59",
   717 => x"78923883",
   718 => x"fff1c40b",
   719 => x"84808080",
   720 => x"b02d5473",
   721 => x"822e8938",
   722 => x"80558480",
   723 => x"809a9504",
   724 => x"83fff1c5",
   725 => x"0b848080",
   726 => x"80b02d70",
   727 => x"83fff5e8",
   728 => x"0cff1170",
   729 => x"83fff5dc",
   730 => x"0c545284",
   731 => x"8080a5f0",
   732 => x"51848080",
   733 => x"81f42d83",
   734 => x"fff1c60b",
   735 => x"84808080",
   736 => x"b02d83ff",
   737 => x"f1c70b84",
   738 => x"808080b0",
   739 => x"2d567605",
   740 => x"75828029",
   741 => x"057083ff",
   742 => x"f5d00c83",
   743 => x"fff1c80b",
   744 => x"84808080",
   745 => x"b02d7083",
   746 => x"fff5c80c",
   747 => x"83fff5e0",
   748 => x"08595758",
   749 => x"76802e81",
   750 => x"ec388853",
   751 => x"848080a4",
   752 => x"b85283ff",
   753 => x"f28a5184",
   754 => x"80809193",
   755 => x"2d785583",
   756 => x"ffe08008",
   757 => x"82bf3883",
   758 => x"fff5e808",
   759 => x"70842b83",
   760 => x"fff5b80c",
   761 => x"7083fff5",
   762 => x"e40c83ff",
   763 => x"f1dd0b84",
   764 => x"808080b0",
   765 => x"2d83fff1",
   766 => x"dc0b8480",
   767 => x"8080b02d",
   768 => x"71828029",
   769 => x"0583fff1",
   770 => x"de0b8480",
   771 => x"8080b02d",
   772 => x"70848080",
   773 => x"291283ff",
   774 => x"f1df0b84",
   775 => x"808080b0",
   776 => x"2d708180",
   777 => x"0a291270",
   778 => x"83fff1b0",
   779 => x"0c83fff5",
   780 => x"c8087129",
   781 => x"83fff5d0",
   782 => x"08057083",
   783 => x"fff5f00c",
   784 => x"83fff1e5",
   785 => x"0b848080",
   786 => x"80b02d83",
   787 => x"fff1e40b",
   788 => x"84808080",
   789 => x"b02d7182",
   790 => x"80290583",
   791 => x"fff1e60b",
   792 => x"84808080",
   793 => x"b02d7084",
   794 => x"80802912",
   795 => x"83fff1e7",
   796 => x"0b848080",
   797 => x"80b02d70",
   798 => x"982b81f0",
   799 => x"0a067205",
   800 => x"7083fff1",
   801 => x"b40cfe11",
   802 => x"7e297705",
   803 => x"83fff5d8",
   804 => x"0c525752",
   805 => x"575d5751",
   806 => x"525f525c",
   807 => x"57575784",
   808 => x"80809a93",
   809 => x"0483fff1",
   810 => x"ca0b8480",
   811 => x"8080b02d",
   812 => x"83fff1c9",
   813 => x"0b848080",
   814 => x"80b02d71",
   815 => x"82802905",
   816 => x"7083fff5",
   817 => x"b80c70a0",
   818 => x"2983ff05",
   819 => x"70892a70",
   820 => x"83fff5e4",
   821 => x"0c83fff1",
   822 => x"cf0b8480",
   823 => x"8080b02d",
   824 => x"83fff1ce",
   825 => x"0b848080",
   826 => x"80b02d71",
   827 => x"82802905",
   828 => x"7083fff1",
   829 => x"b00c7b71",
   830 => x"291e7083",
   831 => x"fff5d80c",
   832 => x"7d83fff1",
   833 => x"b40c7305",
   834 => x"83fff5f0",
   835 => x"0c555e51",
   836 => x"51555581",
   837 => x"557483ff",
   838 => x"e0800c02",
   839 => x"a8050d04",
   840 => x"02ec050d",
   841 => x"7670872c",
   842 => x"7180ff06",
   843 => x"57555383",
   844 => x"fff5e008",
   845 => x"8a387288",
   846 => x"2c7381ff",
   847 => x"06565473",
   848 => x"83fff5cc",
   849 => x"082ebc38",
   850 => x"83fff5d0",
   851 => x"08145284",
   852 => x"8080a694",
   853 => x"51848080",
   854 => x"81f42d83",
   855 => x"fff1b852",
   856 => x"83fff5d0",
   857 => x"08145184",
   858 => x"80808caa",
   859 => x"2d83ffe0",
   860 => x"80085383",
   861 => x"ffe08008",
   862 => x"802e80cf",
   863 => x"387383ff",
   864 => x"f5cc0c83",
   865 => x"fff5e008",
   866 => x"802ea238",
   867 => x"74842983",
   868 => x"fff1b805",
   869 => x"70085253",
   870 => x"8480808d",
   871 => x"e72d83ff",
   872 => x"e08008f0",
   873 => x"0a065584",
   874 => x"80809bc9",
   875 => x"04741083",
   876 => x"fff1b805",
   877 => x"70848080",
   878 => x"809b2d52",
   879 => x"53848080",
   880 => x"8e992d83",
   881 => x"ffe08008",
   882 => x"55745372",
   883 => x"83ffe080",
   884 => x"0c029405",
   885 => x"0d0402c8",
   886 => x"050d7f61",
   887 => x"5f5c8057",
   888 => x"ff0b83ff",
   889 => x"f5cc0c83",
   890 => x"fff1b408",
   891 => x"83fff5d8",
   892 => x"08575883",
   893 => x"fff5e008",
   894 => x"772e8f38",
   895 => x"83fff5e8",
   896 => x"08842b59",
   897 => x"8480809c",
   898 => x"920483ff",
   899 => x"f5e40884",
   900 => x"2b59805a",
   901 => x"79792781",
   902 => x"ea38798f",
   903 => x"06a01858",
   904 => x"5473a438",
   905 => x"75528480",
   906 => x"80a6b451",
   907 => x"84808081",
   908 => x"f42d83ff",
   909 => x"f1b85275",
   910 => x"51811656",
   911 => x"8480808c",
   912 => x"aa2d83ff",
   913 => x"f1b85780",
   914 => x"77848080",
   915 => x"80b02d56",
   916 => x"5474742e",
   917 => x"83388154",
   918 => x"7481e52e",
   919 => x"819c3881",
   920 => x"70750655",
   921 => x"5d73802e",
   922 => x"8190388b",
   923 => x"17848080",
   924 => x"80b02d98",
   925 => x"065b7a81",
   926 => x"81388b53",
   927 => x"7d527651",
   928 => x"84808091",
   929 => x"932d83ff",
   930 => x"e0800880",
   931 => x"ed389c17",
   932 => x"08518480",
   933 => x"808de72d",
   934 => x"83ffe080",
   935 => x"08841d0c",
   936 => x"9a178480",
   937 => x"80809b2d",
   938 => x"51848080",
   939 => x"8e992d83",
   940 => x"ffe08008",
   941 => x"83ffe080",
   942 => x"08881e0c",
   943 => x"83ffe080",
   944 => x"08555583",
   945 => x"fff5e008",
   946 => x"802ea038",
   947 => x"94178480",
   948 => x"80809b2d",
   949 => x"51848080",
   950 => x"8e992d83",
   951 => x"ffe08008",
   952 => x"902b83ff",
   953 => x"f00a0670",
   954 => x"16515473",
   955 => x"881d0c7a",
   956 => x"7c0c7c54",
   957 => x"8480809e",
   958 => x"d504811a",
   959 => x"5a848080",
   960 => x"9c940483",
   961 => x"fff5e008",
   962 => x"802e80c7",
   963 => x"38775184",
   964 => x"80809aa0",
   965 => x"2d83ffe0",
   966 => x"800883ff",
   967 => x"e0800853",
   968 => x"848080a6",
   969 => x"d4525884",
   970 => x"808081f4",
   971 => x"2d7780ff",
   972 => x"fffff806",
   973 => x"547380ff",
   974 => x"fffff82e",
   975 => x"9638fe18",
   976 => x"83fff5e8",
   977 => x"082983ff",
   978 => x"f5f00805",
   979 => x"56848080",
   980 => x"9c920480",
   981 => x"547383ff",
   982 => x"e0800c02",
   983 => x"b8050d04",
   984 => x"02e4050d",
   985 => x"787a7154",
   986 => x"83fff5bc",
   987 => x"53555584",
   988 => x"80809bd6",
   989 => x"2d83ffe0",
   990 => x"800881ff",
   991 => x"06537280",
   992 => x"2e818838",
   993 => x"848080a6",
   994 => x"ec518480",
   995 => x"8084d62d",
   996 => x"83fff5c0",
   997 => x"0883ff05",
   998 => x"892a5780",
   999 => x"70565675",
  1000 => x"77258187",
  1001 => x"3883fff5",
  1002 => x"c408fe05",
  1003 => x"83fff5e8",
  1004 => x"082983ff",
  1005 => x"f5f00811",
  1006 => x"7683fff5",
  1007 => x"dc080605",
  1008 => x"75545253",
  1009 => x"8480808c",
  1010 => x"aa2d83ff",
  1011 => x"e0800880",
  1012 => x"2e80cc38",
  1013 => x"81157083",
  1014 => x"fff5dc08",
  1015 => x"06545572",
  1016 => x"973883ff",
  1017 => x"f5c40851",
  1018 => x"8480809a",
  1019 => x"a02d83ff",
  1020 => x"e0800883",
  1021 => x"fff5c40c",
  1022 => x"84801481",
  1023 => x"17575476",
  1024 => x"7624ffa1",
  1025 => x"38848080",
  1026 => x"a0ab0474",
  1027 => x"52848080",
  1028 => x"a7885184",
  1029 => x"808081f4",
  1030 => x"2d848080",
  1031 => x"a0ad0483",
  1032 => x"ffe08008",
  1033 => x"53848080",
  1034 => x"a0ad0481",
  1035 => x"537283ff",
  1036 => x"e0800c02",
  1037 => x"9c050d04",
  1038 => x"83ffe08c",
  1039 => x"080283ff",
  1040 => x"e08c0cff",
  1041 => x"3d0d800b",
  1042 => x"83ffe08c",
  1043 => x"08fc050c",
  1044 => x"83ffe08c",
  1045 => x"08880508",
  1046 => x"8106ff11",
  1047 => x"70097083",
  1048 => x"ffe08c08",
  1049 => x"8c050806",
  1050 => x"83ffe08c",
  1051 => x"08fc0508",
  1052 => x"1183ffe0",
  1053 => x"8c08fc05",
  1054 => x"0c83ffe0",
  1055 => x"8c088805",
  1056 => x"08812a83",
  1057 => x"ffe08c08",
  1058 => x"88050c83",
  1059 => x"ffe08c08",
  1060 => x"8c050810",
  1061 => x"83ffe08c",
  1062 => x"088c050c",
  1063 => x"51515151",
  1064 => x"83ffe08c",
  1065 => x"08880508",
  1066 => x"802e8438",
  1067 => x"ffa23983",
  1068 => x"ffe08c08",
  1069 => x"fc050870",
  1070 => x"83ffe080",
  1071 => x"0c51833d",
  1072 => x"0d83ffe0",
  1073 => x"8c0c0400",
  1074 => x"00ffffff",
  1075 => x"ff00ffff",
  1076 => x"ffff00ff",
  1077 => x"ffffff00",
  1078 => x"436d645f",
  1079 => x"696e6974",
  1080 => x"0a000000",
  1081 => x"636d645f",
  1082 => x"434d4438",
  1083 => x"20726573",
  1084 => x"706f6e73",
  1085 => x"653a2025",
  1086 => x"640a0000",
  1087 => x"434d4438",
  1088 => x"5f342072",
  1089 => x"6573706f",
  1090 => x"6e73653a",
  1091 => x"2025640a",
  1092 => x"00000000",
  1093 => x"53444843",
  1094 => x"20496e69",
  1095 => x"7469616c",
  1096 => x"697a6174",
  1097 => x"696f6e20",
  1098 => x"6572726f",
  1099 => x"72210a00",
  1100 => x"434d4435",
  1101 => x"38202564",
  1102 => x"0a202000",
  1103 => x"434d4435",
  1104 => x"385f3220",
  1105 => x"25640a20",
  1106 => x"20000000",
  1107 => x"53504920",
  1108 => x"496e6974",
  1109 => x"28290a00",
  1110 => x"52656164",
  1111 => x"20636f6d",
  1112 => x"6d616e64",
  1113 => x"20666169",
  1114 => x"6c656420",
  1115 => x"61742025",
  1116 => x"64202825",
  1117 => x"64290a00",
  1118 => x"496e6974",
  1119 => x"69616c69",
  1120 => x"7a696e67",
  1121 => x"20534420",
  1122 => x"63617264",
  1123 => x"0a000000",
  1124 => x"48756e74",
  1125 => x"696e6720",
  1126 => x"666f7220",
  1127 => x"70617274",
  1128 => x"6974696f",
  1129 => x"6e0a0000",
  1130 => x"4d414e49",
  1131 => x"46455354",
  1132 => x"4d535400",
  1133 => x"50617273",
  1134 => x"696e6720",
  1135 => x"6d616e69",
  1136 => x"66657374",
  1137 => x"0a000000",
  1138 => x"4c6f6164",
  1139 => x"696e6720",
  1140 => x"6d616e69",
  1141 => x"66657374",
  1142 => x"20666169",
  1143 => x"6c65640a",
  1144 => x"00000000",
  1145 => x"52657475",
  1146 => x"726e696e",
  1147 => x"670a0000",
  1148 => x"52656164",
  1149 => x"696e6720",
  1150 => x"4d42520a",
  1151 => x"00000000",
  1152 => x"52656164",
  1153 => x"206f6620",
  1154 => x"4d425220",
  1155 => x"6661696c",
  1156 => x"65640a00",
  1157 => x"4d425220",
  1158 => x"73756363",
  1159 => x"65737366",
  1160 => x"756c6c79",
  1161 => x"20726561",
  1162 => x"640a0000",
  1163 => x"46415431",
  1164 => x"36202020",
  1165 => x"00000000",
  1166 => x"46415433",
  1167 => x"32202020",
  1168 => x"00000000",
  1169 => x"50617274",
  1170 => x"6974696f",
  1171 => x"6e636f75",
  1172 => x"6e742025",
  1173 => x"640a0000",
  1174 => x"4e6f2070",
  1175 => x"61727469",
  1176 => x"74696f6e",
  1177 => x"20736967",
  1178 => x"6e617475",
  1179 => x"72652066",
  1180 => x"6f756e64",
  1181 => x"0a000000",
  1182 => x"52656164",
  1183 => x"696e6720",
  1184 => x"626f6f74",
  1185 => x"20736563",
  1186 => x"746f7220",
  1187 => x"25640a00",
  1188 => x"52656164",
  1189 => x"20626f6f",
  1190 => x"74207365",
  1191 => x"63746f72",
  1192 => x"2066726f",
  1193 => x"6d206669",
  1194 => x"72737420",
  1195 => x"70617274",
  1196 => x"6974696f",
  1197 => x"6e0a0000",
  1198 => x"48756e74",
  1199 => x"696e6720",
  1200 => x"666f7220",
  1201 => x"66696c65",
  1202 => x"73797374",
  1203 => x"656d0a00",
  1204 => x"556e7375",
  1205 => x"70706f72",
  1206 => x"74656420",
  1207 => x"70617274",
  1208 => x"6974696f",
  1209 => x"6e207479",
  1210 => x"7065210d",
  1211 => x"00000000",
  1212 => x"436c7573",
  1213 => x"74657220",
  1214 => x"73697a65",
  1215 => x"3a202564",
  1216 => x"2c20436c",
  1217 => x"75737465",
  1218 => x"72206d61",
  1219 => x"736b2c20",
  1220 => x"25640a00",
  1221 => x"47657443",
  1222 => x"6c757374",
  1223 => x"65722072",
  1224 => x"65616469",
  1225 => x"6e672073",
  1226 => x"6563746f",
  1227 => x"72202564",
  1228 => x"0a000000",
  1229 => x"52656164",
  1230 => x"696e6720",
  1231 => x"64697265",
  1232 => x"63746f72",
  1233 => x"79207365",
  1234 => x"63746f72",
  1235 => x"2025640a",
  1236 => x"00000000",
  1237 => x"47657446",
  1238 => x"41544c69",
  1239 => x"6e6b2072",
  1240 => x"65747572",
  1241 => x"6e656420",
  1242 => x"25640a00",
  1243 => x"4f70656e",
  1244 => x"65642066",
  1245 => x"696c652c",
  1246 => x"206c6f61",
  1247 => x"64696e67",
  1248 => x"2e2e2e0a",
  1249 => x"00000000",
  1250 => x"43616e27",
  1251 => x"74206f70",
  1252 => x"656e2025",
  1253 => x"730a0000",
	others => x"00000000"
);

begin

process (clk)
begin
	if (clk'event and clk = '1') then
		if (from_zpu.memAWriteEnable = '1') and (from_zpu.memBWriteEnable = '1') and (from_zpu.memAAddr=from_zpu.memBAddr) and (from_zpu.memAWrite/=from_zpu.memBWrite) then
			report "write collision" severity failure;
		end if;
	
		if (from_zpu.memAWriteEnable = '1') then
			ram(to_integer(unsigned(from_zpu.memAAddr(maxAddrBitBRAM downto 2)))) := from_zpu.memAWrite;
			to_zpu.memARead <= from_zpu.memAWrite;
		else
			to_zpu.memARead <= ram(to_integer(unsigned(from_zpu.memAAddr(maxAddrBitBRAM downto 2))));
		end if;
	end if;
end process;

process (clk)
begin
	if (clk'event and clk = '1') then
		if (from_zpu.memBWriteEnable = '1') then
			ram(to_integer(unsigned(from_zpu.memBAddr(maxAddrBitBRAM downto 2)))) := from_zpu.memBWrite;
			to_zpu.memBRead <= from_zpu.memBWrite;
		else
			to_zpu.memBRead <= ram(to_integer(unsigned(from_zpu.memBAddr(maxAddrBitBRAM downto 2))));
		end if;
	end if;
end process;


end arch;

