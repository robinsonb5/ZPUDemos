-- ZPU
--
-- Copyright 2004-2008 oharboe - �yvind Harboe - oyvind.harboe@zylin.com
-- Modified by Alastair M. Robinson for the ZPUFlex project.
--
-- The FreeBSD license
-- 
-- Redistribution and use in source and binary forms, with or without
-- modification, are permitted provided that the following conditions
-- are met:
-- 
-- 1. Redistributions of source code must retain the above copyright
--    notice, this list of conditions and the following disclaimer.
-- 2. Redistributions in binary form must reproduce the above
--    copyright notice, this list of conditions and the following
--    disclaimer in the documentation and/or other materials
--    provided with the distribution.
-- 
-- THIS SOFTWARE IS PROVIDED BY THE ZPU PROJECT ``AS IS'' AND ANY
-- EXPRESS OR IMPLIED WARRANTIES, INCLUDING, BUT NOT LIMITED TO,
-- THE IMPLIED WARRANTIES OF MERCHANTABILITY AND FITNESS FOR A
-- PARTICULAR PURPOSE ARE DISCLAIMED. IN NO EVENT SHALL THE
-- ZPU PROJECT OR CONTRIBUTORS BE LIABLE FOR ANY DIRECT,
-- INDIRECT, INCIDENTAL, SPECIAL, EXEMPLARY, OR CONSEQUENTIAL DAMAGES
-- (INCLUDING, BUT NOT LIMITED TO, PROCUREMENT OF SUBSTITUTE GOODS
-- OR SERVICES; LOSS OF USE, DATA, OR PROFITS; OR BUSINESS INTERRUPTION)
-- HOWEVER CAUSED AND ON ANY THEORY OF LIABILITY, WHETHER IN CONTRACT,
-- STRICT LIABILITY, OR TORT (INCLUDING NEGLIGENCE OR OTHERWISE)
-- ARISING IN ANY WAY OUT OF THE USE OF THIS SOFTWARE, EVEN IF
-- ADVISED OF THE POSSIBILITY OF SUCH DAMAGE.
-- 
-- The views and conclusions contained in the software and documentation
-- are those of the authors and should not be interpreted as representing
-- official policies, either expressed or implied, of the ZPU Project.

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;


library work;
use work.zpu_config.all;
use work.zpupkg.all;

entity SDBootstrap_ROM is
generic
	(
		maxAddrBit : integer := maxAddrBitBRAMLimit -- Specify your actual ROM size to save LEs and unnecessary block RAM usage.
	);
port (
	clk : in std_logic;
	areset : in std_logic := '0';
	from_zpu : in ZPU_ToROM;
	to_zpu : out ZPU_FromROM
);
end SDBootstrap_ROM;

architecture arch of SDBootstrap_ROM is

type ram_type is array(natural range 0 to ((2**(maxAddrBit+1))/4)-1) of std_logic_vector(wordSize-1 downto 0);

shared variable ram : ram_type :=
(
     0 => x"0ba08080",
     1 => x"e2040000",
     2 => x"8004a080",
     3 => x"808a0471",
     4 => x"fd060872",
     5 => x"83060981",
     6 => x"05820583",
     7 => x"2b2a83ff",
     8 => x"ff065204",
     9 => x"71fc0608",
    10 => x"72830609",
    11 => x"81058305",
    12 => x"1010102a",
    13 => x"81ff0652",
    14 => x"0471fc06",
    15 => x"080ba080",
    16 => x"9ed07383",
    17 => x"06101005",
    18 => x"08067381",
    19 => x"ff067383",
    20 => x"06098105",
    21 => x"83051010",
    22 => x"102b0772",
    23 => x"fc060c51",
    24 => x"5104a080",
    25 => x"808a0ba0",
    26 => x"808d8204",
    27 => x"0002c405",
    28 => x"0d0280c0",
    29 => x"0583ffe0",
    30 => x"e05b5680",
    31 => x"76708405",
    32 => x"5808715e",
    33 => x"5e577c70",
    34 => x"84055e08",
    35 => x"58805b77",
    36 => x"982a7888",
    37 => x"2b595372",
    38 => x"8838765e",
    39 => x"a0808396",
    40 => x"047b802e",
    41 => x"81ca3880",
    42 => x"5c7280e4",
    43 => x"2e9f3872",
    44 => x"80e4268d",
    45 => x"387280e3",
    46 => x"2e80ee38",
    47 => x"a08082b6",
    48 => x"047280f3",
    49 => x"2e80cc38",
    50 => x"a08082b6",
    51 => x"04758417",
    52 => x"71087e5c",
    53 => x"56575287",
    54 => x"55739c2a",
    55 => x"74842b55",
    56 => x"5271802e",
    57 => x"83388159",
    58 => x"89722589",
    59 => x"38b71252",
    60 => x"a08081f8",
    61 => x"04b01252",
    62 => x"78802e88",
    63 => x"387151a0",
    64 => x"8083a12d",
    65 => x"ff155574",
    66 => x"8025ce38",
    67 => x"8054a080",
    68 => x"82cc0475",
    69 => x"84177108",
    70 => x"70545c57",
    71 => x"52a08083",
    72 => x"c52d7b54",
    73 => x"a08082cc",
    74 => x"04758417",
    75 => x"71085557",
    76 => x"52a08082",
    77 => x"ff04a551",
    78 => x"a08083a1",
    79 => x"2d7251a0",
    80 => x"8083a12d",
    81 => x"821757a0",
    82 => x"80838904",
    83 => x"73ff1555",
    84 => x"52807225",
    85 => x"b4387970",
    86 => x"81055ba0",
    87 => x"8080a42d",
    88 => x"705253a0",
    89 => x"8083a12d",
    90 => x"811757a0",
    91 => x"8082cc04",
    92 => x"72a52e09",
    93 => x"81068838",
    94 => x"815ca080",
    95 => x"83890472",
    96 => x"51a08083",
    97 => x"a12d8117",
    98 => x"57811b5b",
    99 => x"837b25fd",
   100 => x"fe3872fd",
   101 => x"f1387d83",
   102 => x"ffe0800c",
   103 => x"02bc050d",
   104 => x"0402f805",
   105 => x"0d7352c0",
   106 => x"0870882a",
   107 => x"70810651",
   108 => x"51517080",
   109 => x"2ef13871",
   110 => x"c00c7183",
   111 => x"ffe0800c",
   112 => x"0288050d",
   113 => x"0402e805",
   114 => x"0d775574",
   115 => x"70840556",
   116 => x"08538054",
   117 => x"72982a73",
   118 => x"882b5452",
   119 => x"71802ea2",
   120 => x"38c00870",
   121 => x"882a7081",
   122 => x"06515151",
   123 => x"70802ef1",
   124 => x"3871c00c",
   125 => x"81168115",
   126 => x"55568374",
   127 => x"25d63871",
   128 => x"ca387583",
   129 => x"ffe0800c",
   130 => x"0298050d",
   131 => x"0402f405",
   132 => x"0d747671",
   133 => x"81ff06d4",
   134 => x"0c535383",
   135 => x"fff1a008",
   136 => x"85387189",
   137 => x"2b527198",
   138 => x"2ad40c71",
   139 => x"902a7081",
   140 => x"ff06d40c",
   141 => x"5171882a",
   142 => x"7081ff06",
   143 => x"d40c5171",
   144 => x"81ff06d4",
   145 => x"0c72902a",
   146 => x"7081ff06",
   147 => x"d40c51d4",
   148 => x"087081ff",
   149 => x"06515182",
   150 => x"b8bf5270",
   151 => x"81ff2e09",
   152 => x"81069438",
   153 => x"81ff0bd4",
   154 => x"0cd40870",
   155 => x"81ff06ff",
   156 => x"14545151",
   157 => x"71e53870",
   158 => x"83ffe080",
   159 => x"0c028c05",
   160 => x"0d0402fc",
   161 => x"050d81c7",
   162 => x"5181ff0b",
   163 => x"d40cff11",
   164 => x"51708025",
   165 => x"f4380284",
   166 => x"050d0402",
   167 => x"f0050da0",
   168 => x"8085822d",
   169 => x"819c9f53",
   170 => x"805287fc",
   171 => x"80f751a0",
   172 => x"80848d2d",
   173 => x"83ffe080",
   174 => x"085483ff",
   175 => x"e0800881",
   176 => x"2e098106",
   177 => x"ab3881ff",
   178 => x"0bd40c82",
   179 => x"0a52849c",
   180 => x"80e951a0",
   181 => x"80848d2d",
   182 => x"83ffe080",
   183 => x"088d3881",
   184 => x"ff0bd40c",
   185 => x"7353a080",
   186 => x"85f704a0",
   187 => x"8085822d",
   188 => x"ff135372",
   189 => x"ffb23872",
   190 => x"83ffe080",
   191 => x"0c029005",
   192 => x"0d0402f4",
   193 => x"050d81ff",
   194 => x"0bd40ca0",
   195 => x"809ee051",
   196 => x"a08083c5",
   197 => x"2d935380",
   198 => x"5287fc80",
   199 => x"c151a080",
   200 => x"848d2d83",
   201 => x"ffe08008",
   202 => x"8d3881ff",
   203 => x"0bd40c81",
   204 => x"53a08086",
   205 => x"c104a080",
   206 => x"85822dff",
   207 => x"135372d7",
   208 => x"387283ff",
   209 => x"e0800c02",
   210 => x"8c050d04",
   211 => x"02f0050d",
   212 => x"a0808582",
   213 => x"2d83aa52",
   214 => x"849c80c8",
   215 => x"51a08084",
   216 => x"8d2d83ff",
   217 => x"e0800883",
   218 => x"ffe08008",
   219 => x"53a0809e",
   220 => x"ec5254a0",
   221 => x"8080ed2d",
   222 => x"73812e09",
   223 => x"81069038",
   224 => x"d8087083",
   225 => x"ffff0654",
   226 => x"547283aa",
   227 => x"2ea338a0",
   228 => x"8086822d",
   229 => x"a08087aa",
   230 => x"048154a0",
   231 => x"8088df04",
   232 => x"a0809f84",
   233 => x"51a08080",
   234 => x"ed2d8054",
   235 => x"a08088df",
   236 => x"047352a0",
   237 => x"809fa051",
   238 => x"a08080ed",
   239 => x"2d81ff0b",
   240 => x"d40cb153",
   241 => x"a080859b",
   242 => x"2d83ffe0",
   243 => x"8008802e",
   244 => x"80f43880",
   245 => x"5287fc80",
   246 => x"fa51a080",
   247 => x"848d2d83",
   248 => x"ffe08008",
   249 => x"80d03883",
   250 => x"ffe08008",
   251 => x"52a0809f",
   252 => x"b851a080",
   253 => x"80ed2d81",
   254 => x"ff0bd40c",
   255 => x"d40881ff",
   256 => x"067053a0",
   257 => x"809fc452",
   258 => x"54a08080",
   259 => x"ed2d81ff",
   260 => x"0bd40c81",
   261 => x"ff0bd40c",
   262 => x"81ff0bd4",
   263 => x"0c81ff0b",
   264 => x"d40c7386",
   265 => x"2a708106",
   266 => x"70565153",
   267 => x"72802eaf",
   268 => x"38a08087",
   269 => x"990483ff",
   270 => x"e0800852",
   271 => x"a0809fb8",
   272 => x"51a08080",
   273 => x"ed2d7282",
   274 => x"2efed538",
   275 => x"ff135372",
   276 => x"fef238a0",
   277 => x"809fd451",
   278 => x"a08083c5",
   279 => x"2d725473",
   280 => x"83ffe080",
   281 => x"0c029005",
   282 => x"0d0402f4",
   283 => x"050d810b",
   284 => x"83fff1a0",
   285 => x"0cd00870",
   286 => x"8f2a7081",
   287 => x"06515153",
   288 => x"72f33872",
   289 => x"d00ca080",
   290 => x"85822da0",
   291 => x"809fec51",
   292 => x"a08083c5",
   293 => x"2dd00870",
   294 => x"8f2a7081",
   295 => x"06515153",
   296 => x"72f33881",
   297 => x"0bd00c87",
   298 => x"53805284",
   299 => x"d480c051",
   300 => x"a080848d",
   301 => x"2d83ffe0",
   302 => x"8008812e",
   303 => x"09810687",
   304 => x"3883ffe0",
   305 => x"800853a0",
   306 => x"809ffc51",
   307 => x"a08083c5",
   308 => x"2d72822e",
   309 => x"09810692",
   310 => x"38a080a0",
   311 => x"9051a080",
   312 => x"83c52d80",
   313 => x"53a0808a",
   314 => x"da04ff13",
   315 => x"5372ffb9",
   316 => x"38a080a0",
   317 => x"b051a080",
   318 => x"83c52da0",
   319 => x"8086cc2d",
   320 => x"83ffe080",
   321 => x"0883fff1",
   322 => x"a00c83ff",
   323 => x"e0800880",
   324 => x"2e8b38a0",
   325 => x"80a0cc51",
   326 => x"a08083c5",
   327 => x"2da080a0",
   328 => x"e051a080",
   329 => x"83c52d81",
   330 => x"5287fc80",
   331 => x"d051a080",
   332 => x"848d2d81",
   333 => x"ff0bd40c",
   334 => x"d008708f",
   335 => x"2a708106",
   336 => x"51515372",
   337 => x"f33872d0",
   338 => x"0c81ff0b",
   339 => x"d40ca080",
   340 => x"a0f051a0",
   341 => x"8083c52d",
   342 => x"81537283",
   343 => x"ffe0800c",
   344 => x"028c050d",
   345 => x"04800b83",
   346 => x"ffe0800c",
   347 => x"0402e005",
   348 => x"0d797b57",
   349 => x"578058d0",
   350 => x"08708f2a",
   351 => x"70810651",
   352 => x"515473f3",
   353 => x"3882810b",
   354 => x"d00c81ff",
   355 => x"0bd40c76",
   356 => x"5287fc80",
   357 => x"d151a080",
   358 => x"848d2d80",
   359 => x"dbc6df55",
   360 => x"83ffe080",
   361 => x"08802e98",
   362 => x"3883ffe0",
   363 => x"80085376",
   364 => x"52a080a0",
   365 => x"fc51a080",
   366 => x"80ed2da0",
   367 => x"808c8c04",
   368 => x"81ff0bd4",
   369 => x"0cd40870",
   370 => x"81ff0651",
   371 => x"547381fe",
   372 => x"2e098106",
   373 => x"9b3880ff",
   374 => x"55d80876",
   375 => x"70840558",
   376 => x"0cff1555",
   377 => x"748025f1",
   378 => x"388158a0",
   379 => x"808bf604",
   380 => x"ff155574",
   381 => x"cb3881ff",
   382 => x"0bd40cd0",
   383 => x"08708f2a",
   384 => x"70810651",
   385 => x"515473f3",
   386 => x"3873d00c",
   387 => x"7783ffe0",
   388 => x"800c02a0",
   389 => x"050d0402",
   390 => x"f4050d74",
   391 => x"70882a83",
   392 => x"fe800670",
   393 => x"72982a07",
   394 => x"72882b87",
   395 => x"fc808006",
   396 => x"73982b81",
   397 => x"f00a0671",
   398 => x"73070783",
   399 => x"ffe0800c",
   400 => x"56515351",
   401 => x"028c050d",
   402 => x"0402f805",
   403 => x"0d028e05",
   404 => x"a08080a4",
   405 => x"2d74982b",
   406 => x"71902b07",
   407 => x"70902c83",
   408 => x"ffe0800c",
   409 => x"52520288",
   410 => x"050d0402",
   411 => x"f8050d73",
   412 => x"70902b71",
   413 => x"902a0783",
   414 => x"ffe0800c",
   415 => x"52028805",
   416 => x"0d0402ec",
   417 => x"050d800b",
   418 => x"870a0ca0",
   419 => x"80a19c51",
   420 => x"a08083c5",
   421 => x"2da08088",
   422 => x"ea2d83ff",
   423 => x"e0800880",
   424 => x"2e81e638",
   425 => x"a080a1b4",
   426 => x"51a08083",
   427 => x"c52da080",
   428 => x"8fe72d83",
   429 => x"ffe1a052",
   430 => x"a080a1cc",
   431 => x"51a0809b",
   432 => x"f02d83ff",
   433 => x"e0800880",
   434 => x"2e81be38",
   435 => x"83ffe1a0",
   436 => x"0ba080a1",
   437 => x"d85254a0",
   438 => x"8083c52d",
   439 => x"80557370",
   440 => x"810555a0",
   441 => x"8080a42d",
   442 => x"5372a02e",
   443 => x"80de3872",
   444 => x"a32e80fd",
   445 => x"387280c7",
   446 => x"2e098106",
   447 => x"8b38a080",
   448 => x"80882da0",
   449 => x"808ea804",
   450 => x"728a2e09",
   451 => x"81068b38",
   452 => x"a080808a",
   453 => x"2da0808e",
   454 => x"a8047280",
   455 => x"cc2e0981",
   456 => x"06863883",
   457 => x"ffe1a054",
   458 => x"7281df06",
   459 => x"f0057081",
   460 => x"ff065153",
   461 => x"b8732789",
   462 => x"38ef1370",
   463 => x"81ff0651",
   464 => x"5374842b",
   465 => x"730755a0",
   466 => x"808dde04",
   467 => x"72a32ea1",
   468 => x"38737081",
   469 => x"0555a080",
   470 => x"80a42d53",
   471 => x"72a02ef1",
   472 => x"38ff1475",
   473 => x"53705254",
   474 => x"a0809bf0",
   475 => x"2d74870a",
   476 => x"0c737081",
   477 => x"0555a080",
   478 => x"80a42d53",
   479 => x"728a2e09",
   480 => x"8106ee38",
   481 => x"a0808ddc",
   482 => x"04a080a1",
   483 => x"ec51a080",
   484 => x"83c52d80",
   485 => x"0b83ffe0",
   486 => x"800c0294",
   487 => x"050d0402",
   488 => x"e8050d77",
   489 => x"797b5855",
   490 => x"55805372",
   491 => x"7625ab38",
   492 => x"74708105",
   493 => x"56a08080",
   494 => x"a42d7470",
   495 => x"810556a0",
   496 => x"8080a42d",
   497 => x"52527171",
   498 => x"2e883881",
   499 => x"51a0808f",
   500 => x"dc048113",
   501 => x"53a0808f",
   502 => x"ab048051",
   503 => x"7083ffe0",
   504 => x"800c0298",
   505 => x"050d0402",
   506 => x"d8050dff",
   507 => x"0b83fff5",
   508 => x"cc0c800b",
   509 => x"83fff5e0",
   510 => x"0ca080a1",
   511 => x"f851a080",
   512 => x"83c52d83",
   513 => x"fff1b852",
   514 => x"8051a080",
   515 => x"8aed2d83",
   516 => x"ffe08008",
   517 => x"5483ffe0",
   518 => x"80089238",
   519 => x"a080a288",
   520 => x"51a08083",
   521 => x"c52d7355",
   522 => x"a08097cb",
   523 => x"04a080a2",
   524 => x"9c51a080",
   525 => x"83c52d80",
   526 => x"56810b83",
   527 => x"fff1ac0c",
   528 => x"8853a080",
   529 => x"a2b45283",
   530 => x"fff1ee51",
   531 => x"a0808f9f",
   532 => x"2d83ffe0",
   533 => x"8008762e",
   534 => x"0981068b",
   535 => x"3883ffe0",
   536 => x"800883ff",
   537 => x"f1ac0c88",
   538 => x"53a080a2",
   539 => x"c05283ff",
   540 => x"f28a51a0",
   541 => x"808f9f2d",
   542 => x"83ffe080",
   543 => x"088b3883",
   544 => x"ffe08008",
   545 => x"83fff1ac",
   546 => x"0c83fff1",
   547 => x"ac0852a0",
   548 => x"80a2cc51",
   549 => x"a08080ed",
   550 => x"2d83fff1",
   551 => x"ac08802e",
   552 => x"81bb3883",
   553 => x"fff4fe0b",
   554 => x"a08080a4",
   555 => x"2d83fff4",
   556 => x"ff0ba080",
   557 => x"80a42d71",
   558 => x"982b7190",
   559 => x"2b0783ff",
   560 => x"f5800ba0",
   561 => x"8080a42d",
   562 => x"70882b72",
   563 => x"0783fff5",
   564 => x"810ba080",
   565 => x"80a42d71",
   566 => x"0783fff5",
   567 => x"b60ba080",
   568 => x"80a42d83",
   569 => x"fff5b70b",
   570 => x"a08080a4",
   571 => x"2d71882b",
   572 => x"07535f54",
   573 => x"525a5657",
   574 => x"557381ab",
   575 => x"aa2e0981",
   576 => x"06933875",
   577 => x"51a0808c",
   578 => x"972d83ff",
   579 => x"e0800856",
   580 => x"a08092ab",
   581 => x"047382d4",
   582 => x"d52e9038",
   583 => x"a080a2e0",
   584 => x"51a08083",
   585 => x"c52da080",
   586 => x"94a30475",
   587 => x"52a080a3",
   588 => x"8051a080",
   589 => x"80ed2d83",
   590 => x"fff1b852",
   591 => x"7551a080",
   592 => x"8aed2d83",
   593 => x"ffe08008",
   594 => x"5583ffe0",
   595 => x"8008802e",
   596 => x"84f938a0",
   597 => x"80a39851",
   598 => x"a08083c5",
   599 => x"2da080a3",
   600 => x"c051a080",
   601 => x"80ed2d88",
   602 => x"53a080a2",
   603 => x"c05283ff",
   604 => x"f28a51a0",
   605 => x"808f9f2d",
   606 => x"83ffe080",
   607 => x"088d3881",
   608 => x"0b83fff5",
   609 => x"e00ca080",
   610 => x"93b40488",
   611 => x"53a080a2",
   612 => x"b45283ff",
   613 => x"f1ee51a0",
   614 => x"808f9f2d",
   615 => x"83ffe080",
   616 => x"08802e90",
   617 => x"38a080a3",
   618 => x"d851a080",
   619 => x"80ed2da0",
   620 => x"8094a304",
   621 => x"83fff5b6",
   622 => x"0ba08080",
   623 => x"a42d5473",
   624 => x"80d52e09",
   625 => x"810680db",
   626 => x"3883fff5",
   627 => x"b70ba080",
   628 => x"80a42d54",
   629 => x"7381aa2e",
   630 => x"09810680",
   631 => x"c638800b",
   632 => x"83fff1b8",
   633 => x"0ba08080",
   634 => x"a42d5654",
   635 => x"7481e92e",
   636 => x"83388154",
   637 => x"7481eb2e",
   638 => x"8c388055",
   639 => x"73752e09",
   640 => x"810683c7",
   641 => x"3883fff1",
   642 => x"c30ba080",
   643 => x"80a42d55",
   644 => x"74913883",
   645 => x"fff1c40b",
   646 => x"a08080a4",
   647 => x"2d547382",
   648 => x"2e883880",
   649 => x"55a08097",
   650 => x"cb0483ff",
   651 => x"f1c50ba0",
   652 => x"8080a42d",
   653 => x"7083fff5",
   654 => x"e80cff05",
   655 => x"83fff5dc",
   656 => x"0c83fff1",
   657 => x"c60ba080",
   658 => x"80a42d83",
   659 => x"fff1c70b",
   660 => x"a08080a4",
   661 => x"2d587605",
   662 => x"77828029",
   663 => x"057083ff",
   664 => x"f5d00c83",
   665 => x"fff1c80b",
   666 => x"a08080a4",
   667 => x"2d7083ff",
   668 => x"f5c80c83",
   669 => x"fff5e008",
   670 => x"59575876",
   671 => x"802e81df",
   672 => x"388853a0",
   673 => x"80a2c052",
   674 => x"83fff28a",
   675 => x"51a0808f",
   676 => x"9f2d83ff",
   677 => x"e0800882",
   678 => x"b23883ff",
   679 => x"f5e80870",
   680 => x"842b83ff",
   681 => x"f5b80c70",
   682 => x"83fff5e4",
   683 => x"0c83fff1",
   684 => x"dd0ba080",
   685 => x"80a42d83",
   686 => x"fff1dc0b",
   687 => x"a08080a4",
   688 => x"2d718280",
   689 => x"290583ff",
   690 => x"f1de0ba0",
   691 => x"8080a42d",
   692 => x"70848080",
   693 => x"291283ff",
   694 => x"f1df0ba0",
   695 => x"8080a42d",
   696 => x"7081800a",
   697 => x"29127083",
   698 => x"fff1b00c",
   699 => x"83fff5c8",
   700 => x"08712983",
   701 => x"fff5d008",
   702 => x"057083ff",
   703 => x"f5f00c83",
   704 => x"fff1e50b",
   705 => x"a08080a4",
   706 => x"2d83fff1",
   707 => x"e40ba080",
   708 => x"80a42d71",
   709 => x"82802905",
   710 => x"83fff1e6",
   711 => x"0ba08080",
   712 => x"a42d7084",
   713 => x"80802912",
   714 => x"83fff1e7",
   715 => x"0ba08080",
   716 => x"a42d7098",
   717 => x"2b81f00a",
   718 => x"06720570",
   719 => x"83fff1b4",
   720 => x"0cfe117e",
   721 => x"29770583",
   722 => x"fff5d80c",
   723 => x"52595243",
   724 => x"545e5152",
   725 => x"59525d57",
   726 => x"5957a080",
   727 => x"97c90483",
   728 => x"fff1ca0b",
   729 => x"a08080a4",
   730 => x"2d83fff1",
   731 => x"c90ba080",
   732 => x"80a42d71",
   733 => x"82802905",
   734 => x"7083fff5",
   735 => x"b80c70a0",
   736 => x"2983ff05",
   737 => x"70892a70",
   738 => x"83fff5e4",
   739 => x"0c83fff1",
   740 => x"cf0ba080",
   741 => x"80a42d83",
   742 => x"fff1ce0b",
   743 => x"a08080a4",
   744 => x"2d718280",
   745 => x"29057083",
   746 => x"fff1b00c",
   747 => x"7b71291e",
   748 => x"7083fff5",
   749 => x"d80c7d83",
   750 => x"fff1b40c",
   751 => x"730583ff",
   752 => x"f5f00c55",
   753 => x"5e515155",
   754 => x"55815574",
   755 => x"83ffe080",
   756 => x"0c02a805",
   757 => x"0d0402ec",
   758 => x"050d7670",
   759 => x"872c7180",
   760 => x"ff065755",
   761 => x"5383fff5",
   762 => x"e0088a38",
   763 => x"72882c73",
   764 => x"81ff0656",
   765 => x"547383ff",
   766 => x"f5cc082e",
   767 => x"a83883ff",
   768 => x"f1b85283",
   769 => x"fff5d008",
   770 => x"1451a080",
   771 => x"8aed2d83",
   772 => x"ffe08008",
   773 => x"5383ffe0",
   774 => x"8008802e",
   775 => x"80cb3873",
   776 => x"83fff5cc",
   777 => x"0c83fff5",
   778 => x"e008802e",
   779 => x"a0387484",
   780 => x"2983fff1",
   781 => x"b8057008",
   782 => x"5253a080",
   783 => x"8c972d83",
   784 => x"ffe08008",
   785 => x"f00a0655",
   786 => x"a08098e7",
   787 => x"04741083",
   788 => x"fff1b805",
   789 => x"70a08080",
   790 => x"8f2d5253",
   791 => x"a0808cc9",
   792 => x"2d83ffe0",
   793 => x"80085574",
   794 => x"537283ff",
   795 => x"e0800c02",
   796 => x"94050d04",
   797 => x"02cc050d",
   798 => x"7e605e5b",
   799 => x"8056ff0b",
   800 => x"83fff5cc",
   801 => x"0c83fff1",
   802 => x"b40883ff",
   803 => x"f5d80856",
   804 => x"5783fff5",
   805 => x"e008762e",
   806 => x"8e3883ff",
   807 => x"f5e80884",
   808 => x"2b59a080",
   809 => x"99af0483",
   810 => x"fff5e408",
   811 => x"842b5980",
   812 => x"5a797927",
   813 => x"81e13879",
   814 => x"8f06a017",
   815 => x"575473a1",
   816 => x"387452a0",
   817 => x"80a3f851",
   818 => x"a08080ed",
   819 => x"2d83fff1",
   820 => x"b8527451",
   821 => x"811555a0",
   822 => x"808aed2d",
   823 => x"83fff1b8",
   824 => x"568076a0",
   825 => x"8080a42d",
   826 => x"55587378",
   827 => x"2e833881",
   828 => x"587381e5",
   829 => x"2e819838",
   830 => x"81707906",
   831 => x"555c7380",
   832 => x"2e818c38",
   833 => x"8b16a080",
   834 => x"80a42d98",
   835 => x"06587780",
   836 => x"fe388b53",
   837 => x"7c527551",
   838 => x"a0808f9f",
   839 => x"2d83ffe0",
   840 => x"800880eb",
   841 => x"389c1608",
   842 => x"51a0808c",
   843 => x"972d83ff",
   844 => x"e0800884",
   845 => x"1c0c9a16",
   846 => x"a080808f",
   847 => x"2d51a080",
   848 => x"8cc92d83",
   849 => x"ffe08008",
   850 => x"83ffe080",
   851 => x"08555583",
   852 => x"fff5e008",
   853 => x"802e9e38",
   854 => x"9416a080",
   855 => x"808f2d51",
   856 => x"a0808cc9",
   857 => x"2d83ffe0",
   858 => x"8008902b",
   859 => x"83fff00a",
   860 => x"06701651",
   861 => x"5473881c",
   862 => x"0c777b0c",
   863 => x"7c52a080",
   864 => x"a49851a0",
   865 => x"8080ed2d",
   866 => x"7b54a080",
   867 => x"9be50481",
   868 => x"1a5aa080",
   869 => x"99b10483",
   870 => x"fff5e008",
   871 => x"802e80c3",
   872 => x"387651a0",
   873 => x"8097d62d",
   874 => x"83ffe080",
   875 => x"0883ffe0",
   876 => x"800853a0",
   877 => x"80a4ac52",
   878 => x"57a08080",
   879 => x"ed2d7680",
   880 => x"fffffff8",
   881 => x"06547380",
   882 => x"fffffff8",
   883 => x"2e9538fe",
   884 => x"1783fff5",
   885 => x"e8082983",
   886 => x"fff5f008",
   887 => x"0555a080",
   888 => x"99af0480",
   889 => x"547383ff",
   890 => x"e0800c02",
   891 => x"b4050d04",
   892 => x"02e4050d",
   893 => x"787a7154",
   894 => x"83fff5bc",
   895 => x"535555a0",
   896 => x"8098f42d",
   897 => x"83ffe080",
   898 => x"0881ff06",
   899 => x"5372802e",
   900 => x"818338a0",
   901 => x"80a4c451",
   902 => x"a08083c5",
   903 => x"2d83fff5",
   904 => x"c00883ff",
   905 => x"05892a57",
   906 => x"80705656",
   907 => x"75772581",
   908 => x"803883ff",
   909 => x"f5c408fe",
   910 => x"0583fff5",
   911 => x"e8082983",
   912 => x"fff5f008",
   913 => x"117683ff",
   914 => x"f5dc0806",
   915 => x"05755452",
   916 => x"53a0808a",
   917 => x"ed2d83ff",
   918 => x"e0800880",
   919 => x"2e80c738",
   920 => x"81157083",
   921 => x"fff5dc08",
   922 => x"06545572",
   923 => x"963883ff",
   924 => x"f5c40851",
   925 => x"a08097d6",
   926 => x"2d83ffe0",
   927 => x"800883ff",
   928 => x"f5c40c84",
   929 => x"80148117",
   930 => x"57547676",
   931 => x"24ffa338",
   932 => x"a0809db1",
   933 => x"047452a0",
   934 => x"80a4e051",
   935 => x"a08080ed",
   936 => x"2da0809d",
   937 => x"b30483ff",
   938 => x"e0800853",
   939 => x"a0809db3",
   940 => x"04815372",
   941 => x"83ffe080",
   942 => x"0c029c05",
   943 => x"0d0483ff",
   944 => x"e08c0802",
   945 => x"83ffe08c",
   946 => x"0cff3d0d",
   947 => x"800b83ff",
   948 => x"e08c08fc",
   949 => x"050c83ff",
   950 => x"e08c0888",
   951 => x"05088106",
   952 => x"ff117009",
   953 => x"7083ffe0",
   954 => x"8c088c05",
   955 => x"080683ff",
   956 => x"e08c08fc",
   957 => x"05081183",
   958 => x"ffe08c08",
   959 => x"fc050c83",
   960 => x"ffe08c08",
   961 => x"88050881",
   962 => x"2a83ffe0",
   963 => x"8c088805",
   964 => x"0c83ffe0",
   965 => x"8c088c05",
   966 => x"081083ff",
   967 => x"e08c088c",
   968 => x"050c5151",
   969 => x"515183ff",
   970 => x"e08c0888",
   971 => x"0508802e",
   972 => x"8438ffa2",
   973 => x"3983ffe0",
   974 => x"8c08fc05",
   975 => x"087083ff",
   976 => x"e0800c51",
   977 => x"833d0d83",
   978 => x"ffe08c0c",
   979 => x"04000000",
   980 => x"00ffffff",
   981 => x"ff00ffff",
   982 => x"ffff00ff",
   983 => x"ffffff00",
   984 => x"436d645f",
   985 => x"696e6974",
   986 => x"0a000000",
   987 => x"636d645f",
   988 => x"434d4438",
   989 => x"20726573",
   990 => x"706f6e73",
   991 => x"653a2025",
   992 => x"640a0000",
   993 => x"53444843",
   994 => x"20496e69",
   995 => x"7469616c",
   996 => x"697a6174",
   997 => x"696f6e20",
   998 => x"6572726f",
   999 => x"72210a00",
  1000 => x"434d4438",
  1001 => x"5f342072",
  1002 => x"6573706f",
  1003 => x"6e73653a",
  1004 => x"2025640a",
  1005 => x"00000000",
  1006 => x"434d4435",
  1007 => x"38202564",
  1008 => x"0a202000",
  1009 => x"434d4435",
  1010 => x"385f3220",
  1011 => x"25640a20",
  1012 => x"20000000",
  1013 => x"44657465",
  1014 => x"726d696e",
  1015 => x"65642053",
  1016 => x"44484320",
  1017 => x"73746174",
  1018 => x"75730a00",
  1019 => x"41637469",
  1020 => x"76617469",
  1021 => x"6e672043",
  1022 => x"530a0000",
  1023 => x"53656e74",
  1024 => x"20726573",
  1025 => x"65742063",
  1026 => x"6f6d6d61",
  1027 => x"6e640a00",
  1028 => x"53442063",
  1029 => x"61726420",
  1030 => x"696e6974",
  1031 => x"69616c69",
  1032 => x"7a617469",
  1033 => x"6f6e2065",
  1034 => x"72726f72",
  1035 => x"210a0000",
  1036 => x"43617264",
  1037 => x"20726573",
  1038 => x"706f6e64",
  1039 => x"65642074",
  1040 => x"6f207265",
  1041 => x"7365740a",
  1042 => x"00000000",
  1043 => x"53444843",
  1044 => x"20636172",
  1045 => x"64206465",
  1046 => x"74656374",
  1047 => x"65640a00",
  1048 => x"53656e64",
  1049 => x"696e6720",
  1050 => x"636d6431",
  1051 => x"360a0000",
  1052 => x"496e6974",
  1053 => x"20646f6e",
  1054 => x"650a0000",
  1055 => x"52656164",
  1056 => x"20636f6d",
  1057 => x"6d616e64",
  1058 => x"20666169",
  1059 => x"6c656420",
  1060 => x"61742025",
  1061 => x"64202825",
  1062 => x"64290a00",
  1063 => x"496e6974",
  1064 => x"69616c69",
  1065 => x"7a696e67",
  1066 => x"20534420",
  1067 => x"63617264",
  1068 => x"0a000000",
  1069 => x"48756e74",
  1070 => x"696e6720",
  1071 => x"666f7220",
  1072 => x"70617274",
  1073 => x"6974696f",
  1074 => x"6e0a0000",
  1075 => x"4d414e49",
  1076 => x"46455354",
  1077 => x"4d535400",
  1078 => x"50617273",
  1079 => x"696e6720",
  1080 => x"6d616e69",
  1081 => x"66657374",
  1082 => x"0a000000",
  1083 => x"52657475",
  1084 => x"726e696e",
  1085 => x"670a0000",
  1086 => x"52656164",
  1087 => x"696e6720",
  1088 => x"4d42520a",
  1089 => x"00000000",
  1090 => x"52656164",
  1091 => x"206f6620",
  1092 => x"4d425220",
  1093 => x"6661696c",
  1094 => x"65640a00",
  1095 => x"4d425220",
  1096 => x"73756363",
  1097 => x"65737366",
  1098 => x"756c6c79",
  1099 => x"20726561",
  1100 => x"640a0000",
  1101 => x"46415431",
  1102 => x"36202020",
  1103 => x"00000000",
  1104 => x"46415433",
  1105 => x"32202020",
  1106 => x"00000000",
  1107 => x"50617274",
  1108 => x"6974696f",
  1109 => x"6e636f75",
  1110 => x"6e742025",
  1111 => x"640a0000",
  1112 => x"4e6f2070",
  1113 => x"61727469",
  1114 => x"74696f6e",
  1115 => x"20736967",
  1116 => x"6e617475",
  1117 => x"72652066",
  1118 => x"6f756e64",
  1119 => x"0a000000",
  1120 => x"52656164",
  1121 => x"696e6720",
  1122 => x"626f6f74",
  1123 => x"20736563",
  1124 => x"746f7220",
  1125 => x"25640a00",
  1126 => x"52656164",
  1127 => x"20626f6f",
  1128 => x"74207365",
  1129 => x"63746f72",
  1130 => x"2066726f",
  1131 => x"6d206669",
  1132 => x"72737420",
  1133 => x"70617274",
  1134 => x"6974696f",
  1135 => x"6e0a0000",
  1136 => x"48756e74",
  1137 => x"696e6720",
  1138 => x"666f7220",
  1139 => x"66696c65",
  1140 => x"73797374",
  1141 => x"656d0a00",
  1142 => x"556e7375",
  1143 => x"70706f72",
  1144 => x"74656420",
  1145 => x"70617274",
  1146 => x"6974696f",
  1147 => x"6e207479",
  1148 => x"7065210d",
  1149 => x"00000000",
  1150 => x"52656164",
  1151 => x"696e6720",
  1152 => x"64697265",
  1153 => x"63746f72",
  1154 => x"79207365",
  1155 => x"63746f72",
  1156 => x"2025640a",
  1157 => x"00000000",
  1158 => x"66696c65",
  1159 => x"20222573",
  1160 => x"2220666f",
  1161 => x"756e640d",
  1162 => x"00000000",
  1163 => x"47657446",
  1164 => x"41544c69",
  1165 => x"6e6b2072",
  1166 => x"65747572",
  1167 => x"6e656420",
  1168 => x"25640a00",
  1169 => x"4f70656e",
  1170 => x"65642066",
  1171 => x"696c652c",
  1172 => x"206c6f61",
  1173 => x"64696e67",
  1174 => x"2e2e2e0a",
  1175 => x"00000000",
  1176 => x"43616e27",
  1177 => x"74206f70",
  1178 => x"656e2025",
  1179 => x"730a0000",
	others => x"00000000"
);

begin

process (clk)
begin
	if (clk'event and clk = '1') then
		if (from_zpu.memAWriteEnable = '1') and (from_zpu.memBWriteEnable = '1') and (from_zpu.memAAddr=from_zpu.memBAddr) and (from_zpu.memAWrite/=from_zpu.memBWrite) then
			report "write collision" severity failure;
		end if;
	
		if (from_zpu.memAWriteEnable = '1') then
			ram(to_integer(unsigned(from_zpu.memAAddr(maxAddrBit downto 2)))) := from_zpu.memAWrite;
			to_zpu.memARead <= from_zpu.memAWrite;
		else
			to_zpu.memARead <= ram(to_integer(unsigned(from_zpu.memAAddr(maxAddrBit downto 2))));
		end if;
	end if;
end process;

process (clk)
begin
	if (clk'event and clk = '1') then
		if (from_zpu.memBWriteEnable = '1') then
			ram(to_integer(unsigned(from_zpu.memBAddr(maxAddrBit downto 2)))) := from_zpu.memBWrite;
			to_zpu.memBRead <= from_zpu.memBWrite;
		else
			to_zpu.memBRead <= ram(to_integer(unsigned(from_zpu.memBAddr(maxAddrBit downto 2))));
		end if;
	end if;
end process;


end arch;

