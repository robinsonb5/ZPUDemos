-- ZPU
--
-- Copyright 2004-2008 oharboe - �yvind Harboe - oyvind.harboe@zylin.com
-- Modified by Alastair M. Robinson for the ZPUFlex project.
--
-- The FreeBSD license
-- 
-- Redistribution and use in source and binary forms, with or without
-- modification, are permitted provided that the following conditions
-- are met:
-- 
-- 1. Redistributions of source code must retain the above copyright
--    notice, this list of conditions and the following disclaimer.
-- 2. Redistributions in binary form must reproduce the above
--    copyright notice, this list of conditions and the following
--    disclaimer in the documentation and/or other materials
--    provided with the distribution.
-- 
-- THIS SOFTWARE IS PROVIDED BY THE ZPU PROJECT ``AS IS'' AND ANY
-- EXPRESS OR IMPLIED WARRANTIES, INCLUDING, BUT NOT LIMITED TO,
-- THE IMPLIED WARRANTIES OF MERCHANTABILITY AND FITNESS FOR A
-- PARTICULAR PURPOSE ARE DISCLAIMED. IN NO EVENT SHALL THE
-- ZPU PROJECT OR CONTRIBUTORS BE LIABLE FOR ANY DIRECT,
-- INDIRECT, INCIDENTAL, SPECIAL, EXEMPLARY, OR CONSEQUENTIAL DAMAGES
-- (INCLUDING, BUT NOT LIMITED TO, PROCUREMENT OF SUBSTITUTE GOODS
-- OR SERVICES; LOSS OF USE, DATA, OR PROFITS; OR BUSINESS INTERRUPTION)
-- HOWEVER CAUSED AND ON ANY THEORY OF LIABILITY, WHETHER IN CONTRACT,
-- STRICT LIABILITY, OR TORT (INCLUDING NEGLIGENCE OR OTHERWISE)
-- ARISING IN ANY WAY OUT OF THE USE OF THIS SOFTWARE, EVEN IF
-- ADVISED OF THE POSSIBILITY OF SUCH DAMAGE.
-- 
-- The views and conclusions contained in the software and documentation
-- are those of the authors and should not be interpreted as representing
-- official policies, either expressed or implied, of the ZPU Project.

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;


library work;
use work.zpupkg.all;

entity VGATest_ROM is
generic
	(
		maxAddrBitBRAM : integer := maxAddrBitBRAMLimit -- Specify your actual ROM size to save LEs and unnecessary block RAM usage.
	);
port (
	clk : in std_logic;
	areset : in std_logic := '0';
	from_zpu : in ZPU_ToROM;
	to_zpu : out ZPU_FromROM
);
end VGATest_ROM;

architecture arch of VGATest_ROM is

type ram_type is array(natural range 0 to ((2**(maxAddrBitBRAM+1))/4)-1) of std_logic_vector(wordSize-1 downto 0);

shared variable ram : ram_type :=
(
     0 => x"84808080",
     1 => x"8c0b8480",
     2 => x"8081e004",
     3 => x"00848080",
     4 => x"808c04ff",
     5 => x"0d800404",
     6 => x"40000017",
     7 => x"00000000",
     8 => x"84808098",
     9 => x"c8088480",
    10 => x"8098cc08",
    11 => x"84808098",
    12 => x"d0088480",
    13 => x"80809808",
    14 => x"2d848080",
    15 => x"98d00c84",
    16 => x"808098cc",
    17 => x"0c848080",
    18 => x"98c80c04",
    19 => x"00000000",
    20 => x"00000000",
    21 => x"00000000",
    22 => x"00000000",
    23 => x"00000000",
    24 => x"71fd0608",
    25 => x"72830609",
    26 => x"81058205",
    27 => x"832b2a83",
    28 => x"ffff0652",
    29 => x"0471fc06",
    30 => x"08728306",
    31 => x"09810583",
    32 => x"05101010",
    33 => x"2a81ff06",
    34 => x"520471fd",
    35 => x"060883ff",
    36 => x"ff738306",
    37 => x"09810582",
    38 => x"05832b2b",
    39 => x"09067383",
    40 => x"ffff0673",
    41 => x"83060981",
    42 => x"05820583",
    43 => x"2b0b2b07",
    44 => x"72fc060c",
    45 => x"51510471",
    46 => x"fc060884",
    47 => x"808092bc",
    48 => x"73830610",
    49 => x"10050806",
    50 => x"7381ff06",
    51 => x"73830609",
    52 => x"81058305",
    53 => x"1010102b",
    54 => x"0772fc06",
    55 => x"0c515104",
    56 => x"84808098",
    57 => x"c8708480",
    58 => x"8099e827",
    59 => x"8e388071",
    60 => x"70840553",
    61 => x"0c848080",
    62 => x"81e50484",
    63 => x"8080808c",
    64 => x"51848080",
    65 => x"86cb0402",
    66 => x"c0050d02",
    67 => x"80c4055b",
    68 => x"80707c70",
    69 => x"84055e08",
    70 => x"725f5f5f",
    71 => x"5a7c7084",
    72 => x"055e0857",
    73 => x"80597698",
    74 => x"2a77882b",
    75 => x"58557480",
    76 => x"2e82e738",
    77 => x"7b802e80",
    78 => x"d338805c",
    79 => x"7480e42e",
    80 => x"81d83874",
    81 => x"80f82e81",
    82 => x"d1387480",
    83 => x"e42e81dc",
    84 => x"387480e4",
    85 => x"2680f138",
    86 => x"7480e32e",
    87 => x"80c838a5",
    88 => x"51848080",
    89 => x"85db2d74",
    90 => x"51848080",
    91 => x"85db2d82",
    92 => x"1a811a5a",
    93 => x"5a837925",
    94 => x"ffac3874",
    95 => x"ff9f387e",
    96 => x"84808098",
    97 => x"c80c0280",
    98 => x"c0050d04",
    99 => x"74a52e09",
   100 => x"81069b38",
   101 => x"810b811a",
   102 => x"5a5c8379",
   103 => x"25ff8738",
   104 => x"84808082",
   105 => x"fb047a84",
   106 => x"1c710857",
   107 => x"5c547451",
   108 => x"84808085",
   109 => x"db2d811a",
   110 => x"811a5a5a",
   111 => x"837925fe",
   112 => x"e5388480",
   113 => x"8082fb04",
   114 => x"7480f32e",
   115 => x"81d93874",
   116 => x"80f82e09",
   117 => x"8106ff87",
   118 => x"387d5380",
   119 => x"587d782e",
   120 => x"81e23887",
   121 => x"56729c2a",
   122 => x"73842b54",
   123 => x"5271802e",
   124 => x"83388158",
   125 => x"b7125471",
   126 => x"89248438",
   127 => x"b0125477",
   128 => x"80ea38ff",
   129 => x"16567580",
   130 => x"25db3881",
   131 => x"19598379",
   132 => x"25fe9338",
   133 => x"84808082",
   134 => x"fb047a84",
   135 => x"1c710840",
   136 => x"5c527480",
   137 => x"e42e0981",
   138 => x"06fea638",
   139 => x"7d538058",
   140 => x"7d782e81",
   141 => x"8f388756",
   142 => x"729c2a73",
   143 => x"842b5452",
   144 => x"71802e83",
   145 => x"388158b7",
   146 => x"12547189",
   147 => x"248438b0",
   148 => x"125477af",
   149 => x"38ff1656",
   150 => x"758025dc",
   151 => x"38811959",
   152 => x"837925fd",
   153 => x"c1388480",
   154 => x"8082fb04",
   155 => x"73518480",
   156 => x"8085db2d",
   157 => x"ff165675",
   158 => x"8025fee9",
   159 => x"38848080",
   160 => x"848b0473",
   161 => x"51848080",
   162 => x"85db2dff",
   163 => x"16567580",
   164 => x"25ffa538",
   165 => x"84808084",
   166 => x"dd047984",
   167 => x"808098c8",
   168 => x"0c0280c0",
   169 => x"050d047a",
   170 => x"841c7108",
   171 => x"535c5384",
   172 => x"80808680",
   173 => x"2d811959",
   174 => x"837925fc",
   175 => x"e9388480",
   176 => x"8082fb04",
   177 => x"b0518480",
   178 => x"8085db2d",
   179 => x"81195983",
   180 => x"7925fcd2",
   181 => x"38848080",
   182 => x"82fb0402",
   183 => x"f8050d73",
   184 => x"52c00870",
   185 => x"882a7081",
   186 => x"06515151",
   187 => x"70802ef1",
   188 => x"3871c00c",
   189 => x"71848080",
   190 => x"98c80c02",
   191 => x"88050d04",
   192 => x"02e8050d",
   193 => x"80785755",
   194 => x"75708405",
   195 => x"57085380",
   196 => x"5472982a",
   197 => x"73882b54",
   198 => x"5271802e",
   199 => x"a238c008",
   200 => x"70882a70",
   201 => x"81065151",
   202 => x"5170802e",
   203 => x"f13871c0",
   204 => x"0c811581",
   205 => x"15555583",
   206 => x"7425d638",
   207 => x"71ca3874",
   208 => x"84808098",
   209 => x"c80c0298",
   210 => x"050d0402",
   211 => x"e8050d80",
   212 => x"56848080",
   213 => x"0bfc800c",
   214 => x"81167057",
   215 => x"52848080",
   216 => x"54805584",
   217 => x"fe538112",
   218 => x"7083ffff",
   219 => x"06707670",
   220 => x"8405580c",
   221 => x"fe155551",
   222 => x"52728025",
   223 => x"e9388115",
   224 => x"5583df75",
   225 => x"25dd3880",
   226 => x"51848080",
   227 => x"8efa2d84",
   228 => x"808086d8",
   229 => x"0402f405",
   230 => x"0d747652",
   231 => x"53807125",
   232 => x"90387052",
   233 => x"72708405",
   234 => x"5408ff13",
   235 => x"535171f4",
   236 => x"38028c05",
   237 => x"0d0402d4",
   238 => x"050d7c7e",
   239 => x"5c58810b",
   240 => x"84808092",
   241 => x"cc585a83",
   242 => x"59760878",
   243 => x"0c770877",
   244 => x"08565473",
   245 => x"752e9438",
   246 => x"77085374",
   247 => x"52848080",
   248 => x"92dc5184",
   249 => x"80808287",
   250 => x"2d805a77",
   251 => x"56807b25",
   252 => x"90387a55",
   253 => x"75708405",
   254 => x"5708ff16",
   255 => x"565474f4",
   256 => x"38770877",
   257 => x"08565675",
   258 => x"752e9438",
   259 => x"77085374",
   260 => x"52848080",
   261 => x"939c5184",
   262 => x"80808287",
   263 => x"2d805aff",
   264 => x"19841858",
   265 => x"59788025",
   266 => x"ff9f3879",
   267 => x"84808098",
   268 => x"c80c02ac",
   269 => x"050d0402",
   270 => x"e4050d78",
   271 => x"7a555681",
   272 => x"5785aad5",
   273 => x"aad5760c",
   274 => x"fad5aad5",
   275 => x"aa0b8c17",
   276 => x"0ccc7684",
   277 => x"808081b7",
   278 => x"2db30b8f",
   279 => x"17848080",
   280 => x"81b72d75",
   281 => x"085372fc",
   282 => x"e2d5aad5",
   283 => x"2e923875",
   284 => x"08528480",
   285 => x"8093dc51",
   286 => x"84808082",
   287 => x"872d8057",
   288 => x"8c160855",
   289 => x"74fad5aa",
   290 => x"d4b32e93",
   291 => x"388c1608",
   292 => x"52848080",
   293 => x"94985184",
   294 => x"80808287",
   295 => x"2d805775",
   296 => x"55807425",
   297 => x"8e387470",
   298 => x"84055608",
   299 => x"ff155553",
   300 => x"73f43875",
   301 => x"085473fc",
   302 => x"e2d5aad5",
   303 => x"2e923875",
   304 => x"08528480",
   305 => x"8094d451",
   306 => x"84808082",
   307 => x"872d8057",
   308 => x"8c160853",
   309 => x"72fad5aa",
   310 => x"d4b32e93",
   311 => x"388c1608",
   312 => x"52848080",
   313 => x"95905184",
   314 => x"80808287",
   315 => x"2d805776",
   316 => x"84808098",
   317 => x"c80c029c",
   318 => x"050d0402",
   319 => x"c4050d60",
   320 => x"5c806290",
   321 => x"808029ff",
   322 => x"05848080",
   323 => x"95cc535a",
   324 => x"5b848080",
   325 => x"82872d80",
   326 => x"e1b35782",
   327 => x"5fae5184",
   328 => x"808085db",
   329 => x"2d761070",
   330 => x"962a8106",
   331 => x"56577480",
   332 => x"2e853876",
   333 => x"81075776",
   334 => x"952a8106",
   335 => x"5877802e",
   336 => x"85387681",
   337 => x"32577977",
   338 => x"07790677",
   339 => x"5f5a8fff",
   340 => x"ff587679",
   341 => x"06707b32",
   342 => x"822b7d11",
   343 => x"5157760c",
   344 => x"76107096",
   345 => x"2a810656",
   346 => x"5774802e",
   347 => x"85387681",
   348 => x"07577695",
   349 => x"2a810655",
   350 => x"74802e85",
   351 => x"38768132",
   352 => x"57ff1858",
   353 => x"778025ca",
   354 => x"387d578f",
   355 => x"ffff5876",
   356 => x"7906707b",
   357 => x"32822b7d",
   358 => x"05700857",
   359 => x"5f567476",
   360 => x"2e80ea38",
   361 => x"807b5384",
   362 => x"808095dc",
   363 => x"525d8480",
   364 => x"8082872d",
   365 => x"74547553",
   366 => x"75528480",
   367 => x"8095f051",
   368 => x"84808082",
   369 => x"872d7c5b",
   370 => x"76107096",
   371 => x"2a810657",
   372 => x"5775802e",
   373 => x"85387681",
   374 => x"07577695",
   375 => x"2a810655",
   376 => x"74802e85",
   377 => x"38768132",
   378 => x"57ff1858",
   379 => x"778025ff",
   380 => x"9e38ff1f",
   381 => x"5f7efea5",
   382 => x"388a5184",
   383 => x"808085db",
   384 => x"2d7c8480",
   385 => x"8098c80c",
   386 => x"02bc050d",
   387 => x"04811b5b",
   388 => x"8480808b",
   389 => x"c80402cc",
   390 => x"050d7e60",
   391 => x"5e58815a",
   392 => x"805b80c0",
   393 => x"7a585c85",
   394 => x"ada989bb",
   395 => x"780c7959",
   396 => x"81569755",
   397 => x"76760782",
   398 => x"2b781151",
   399 => x"5485ada9",
   400 => x"89bb740c",
   401 => x"7510ff16",
   402 => x"56567480",
   403 => x"25e63876",
   404 => x"10811a5a",
   405 => x"57987925",
   406 => x"d7387756",
   407 => x"807d2590",
   408 => x"387c5575",
   409 => x"70840557",
   410 => x"08ff1656",
   411 => x"5474f438",
   412 => x"8157ff87",
   413 => x"87a5c378",
   414 => x"0c975976",
   415 => x"822b7811",
   416 => x"70085f56",
   417 => x"567cff87",
   418 => x"87a5c32e",
   419 => x"80cc3874",
   420 => x"08547385",
   421 => x"ada989bb",
   422 => x"2e943880",
   423 => x"75085476",
   424 => x"53848080",
   425 => x"9698525a",
   426 => x"84808082",
   427 => x"872d7610",
   428 => x"ff1a5a57",
   429 => x"788025c3",
   430 => x"387a822b",
   431 => x"5675b138",
   432 => x"7b528480",
   433 => x"8096b851",
   434 => x"84808082",
   435 => x"872d7b84",
   436 => x"808098c8",
   437 => x"0c02b405",
   438 => x"0d047a77",
   439 => x"077710ff",
   440 => x"1b5b585b",
   441 => x"788025ff",
   442 => x"92388480",
   443 => x"808db904",
   444 => x"75528480",
   445 => x"8096f451",
   446 => x"84808082",
   447 => x"872d7599",
   448 => x"2a813281",
   449 => x"06700981",
   450 => x"05710770",
   451 => x"09709f2c",
   452 => x"7d067910",
   453 => x"9ffffffc",
   454 => x"0660812a",
   455 => x"415a5d57",
   456 => x"585975da",
   457 => x"38790981",
   458 => x"05707b07",
   459 => x"9f2a5556",
   460 => x"7bbf2684",
   461 => x"38739d38",
   462 => x"81705384",
   463 => x"808096b8",
   464 => x"525c8480",
   465 => x"8082872d",
   466 => x"7b848080",
   467 => x"98c80c02",
   468 => x"b4050d04",
   469 => x"84808097",
   470 => x"8c518480",
   471 => x"8082872d",
   472 => x"7b528480",
   473 => x"8096b851",
   474 => x"84808082",
   475 => x"872d7b84",
   476 => x"808098c8",
   477 => x"0c02b405",
   478 => x"0d0402d4",
   479 => x"050d7c57",
   480 => x"81708480",
   481 => x"8092cc5b",
   482 => x"595b835a",
   483 => x"7808770c",
   484 => x"76087908",
   485 => x"56547375",
   486 => x"2e943876",
   487 => x"08537452",
   488 => x"84808092",
   489 => x"dc518480",
   490 => x"8082872d",
   491 => x"80587656",
   492 => x"9fff5575",
   493 => x"70840557",
   494 => x"08ff1656",
   495 => x"54748025",
   496 => x"f2387608",
   497 => x"79085656",
   498 => x"75752e94",
   499 => x"38760853",
   500 => x"74528480",
   501 => x"80939c51",
   502 => x"84808082",
   503 => x"872d8058",
   504 => x"ff1a841a",
   505 => x"5a5a7980",
   506 => x"25ffa138",
   507 => x"7781fd38",
   508 => x"775b8158",
   509 => x"85aad5aa",
   510 => x"d5770cfa",
   511 => x"d5aad5aa",
   512 => x"0b8c180c",
   513 => x"cc778480",
   514 => x"8081b72d",
   515 => x"b30b8f18",
   516 => x"84808081",
   517 => x"b72d7608",
   518 => x"5574fce2",
   519 => x"d5aad52e",
   520 => x"92387608",
   521 => x"52848080",
   522 => x"93dc5184",
   523 => x"80808287",
   524 => x"2d80588c",
   525 => x"17085978",
   526 => x"fad5aad4",
   527 => x"b32e9338",
   528 => x"8c170852",
   529 => x"84808094",
   530 => x"98518480",
   531 => x"8082872d",
   532 => x"80587656",
   533 => x"9fff5575",
   534 => x"70840557",
   535 => x"08ff1656",
   536 => x"54748025",
   537 => x"f2387608",
   538 => x"5a79fce2",
   539 => x"d5aad52e",
   540 => x"92387608",
   541 => x"52848080",
   542 => x"94d45184",
   543 => x"80808287",
   544 => x"2d80588c",
   545 => x"17085473",
   546 => x"fad5aad4",
   547 => x"b32e80ee",
   548 => x"388c1708",
   549 => x"52848080",
   550 => x"95905184",
   551 => x"80808287",
   552 => x"2d805877",
   553 => x"5ba08052",
   554 => x"76518480",
   555 => x"808c962d",
   556 => x"84808098",
   557 => x"c8085484",
   558 => x"808098c8",
   559 => x"0880e938",
   560 => x"84808098",
   561 => x"c8085b73",
   562 => x"52765184",
   563 => x"808089fb",
   564 => x"2d848080",
   565 => x"98c808be",
   566 => x"38848080",
   567 => x"98c8085b",
   568 => x"7a848080",
   569 => x"98c80c02",
   570 => x"ac050d04",
   571 => x"84808097",
   572 => x"d8518480",
   573 => x"8082872d",
   574 => x"8480808f",
   575 => x"f2047780",
   576 => x"2effa038",
   577 => x"84808097",
   578 => x"fc518480",
   579 => x"8082872d",
   580 => x"84808091",
   581 => x"a5048480",
   582 => x"80989851",
   583 => x"84808082",
   584 => x"872d8480",
   585 => x"8091e004",
   586 => x"84808098",
   587 => x"b0518480",
   588 => x"8082872d",
   589 => x"84808091",
   590 => x"c7040000",
   591 => x"00ffffff",
   592 => x"ff00ffff",
   593 => x"ffff00ff",
   594 => x"ffffff00",
   595 => x"00000000",
   596 => x"55555555",
   597 => x"aaaaaaaa",
   598 => x"ffffffff",
   599 => x"53616e69",
   600 => x"74792063",
   601 => x"6865636b",
   602 => x"20666169",
   603 => x"6c656420",
   604 => x"28626566",
   605 => x"6f726520",
   606 => x"63616368",
   607 => x"65207265",
   608 => x"66726573",
   609 => x"6829206f",
   610 => x"6e203078",
   611 => x"25642028",
   612 => x"676f7420",
   613 => x"30782564",
   614 => x"290a0000",
   615 => x"53616e69",
   616 => x"74792063",
   617 => x"6865636b",
   618 => x"20666169",
   619 => x"6c656420",
   620 => x"28616674",
   621 => x"65722063",
   622 => x"61636865",
   623 => x"20726566",
   624 => x"72657368",
   625 => x"29206f6e",
   626 => x"20307825",
   627 => x"64202867",
   628 => x"6f742030",
   629 => x"78256429",
   630 => x"0a000000",
   631 => x"42797465",
   632 => x"20636865",
   633 => x"636b2066",
   634 => x"61696c65",
   635 => x"64202862",
   636 => x"65666f72",
   637 => x"65206361",
   638 => x"63686520",
   639 => x"72656672",
   640 => x"65736829",
   641 => x"20617420",
   642 => x"30202867",
   643 => x"6f742030",
   644 => x"78256429",
   645 => x"0a000000",
   646 => x"42797465",
   647 => x"20636865",
   648 => x"636b2066",
   649 => x"61696c65",
   650 => x"64202862",
   651 => x"65666f72",
   652 => x"65206361",
   653 => x"63686520",
   654 => x"72656672",
   655 => x"65736829",
   656 => x"20617420",
   657 => x"33202867",
   658 => x"6f742030",
   659 => x"78256429",
   660 => x"0a000000",
   661 => x"42797465",
   662 => x"20636865",
   663 => x"636b2066",
   664 => x"61696c65",
   665 => x"64202861",
   666 => x"66746572",
   667 => x"20636163",
   668 => x"68652072",
   669 => x"65667265",
   670 => x"73682920",
   671 => x"61742030",
   672 => x"2028676f",
   673 => x"74203078",
   674 => x"2564290a",
   675 => x"00000000",
   676 => x"42797465",
   677 => x"20636865",
   678 => x"636b2066",
   679 => x"61696c65",
   680 => x"64202861",
   681 => x"66746572",
   682 => x"20636163",
   683 => x"68652072",
   684 => x"65667265",
   685 => x"73682920",
   686 => x"61742033",
   687 => x"2028676f",
   688 => x"74203078",
   689 => x"2564290a",
   690 => x"00000000",
   691 => x"43686563",
   692 => x"6b696e67",
   693 => x"206d656d",
   694 => x"6f727900",
   695 => x"30782564",
   696 => x"20676f6f",
   697 => x"64207265",
   698 => x"6164732c",
   699 => x"20000000",
   700 => x"4572726f",
   701 => x"72206174",
   702 => x"20307825",
   703 => x"642c2065",
   704 => x"78706563",
   705 => x"74656420",
   706 => x"30782564",
   707 => x"2c20676f",
   708 => x"74203078",
   709 => x"25640a00",
   710 => x"42616420",
   711 => x"64617461",
   712 => x"20666f75",
   713 => x"6e642061",
   714 => x"74203078",
   715 => x"25642028",
   716 => x"30782564",
   717 => x"290a0000",
   718 => x"53445241",
   719 => x"4d207369",
   720 => x"7a652028",
   721 => x"61737375",
   722 => x"6d696e67",
   723 => x"206e6f20",
   724 => x"61646472",
   725 => x"65737320",
   726 => x"6661756c",
   727 => x"74732920",
   728 => x"69732030",
   729 => x"78256420",
   730 => x"6d656761",
   731 => x"62797465",
   732 => x"730a0000",
   733 => x"416c6961",
   734 => x"73657320",
   735 => x"666f756e",
   736 => x"64206174",
   737 => x"20307825",
   738 => x"640a0000",
   739 => x"28416c69",
   740 => x"61736573",
   741 => x"2070726f",
   742 => x"6261626c",
   743 => x"79207369",
   744 => x"6d706c79",
   745 => x"20696e64",
   746 => x"69636174",
   747 => x"65207468",
   748 => x"61742052",
   749 => x"414d0a69",
   750 => x"7320736d",
   751 => x"616c6c65",
   752 => x"72207468",
   753 => x"616e2036",
   754 => x"34206d65",
   755 => x"67616279",
   756 => x"74657329",
   757 => x"0a000000",
   758 => x"46697273",
   759 => x"74207374",
   760 => x"61676520",
   761 => x"73616e69",
   762 => x"74792063",
   763 => x"6865636b",
   764 => x"20706173",
   765 => x"7365642e",
   766 => x"0a000000",
   767 => x"42797465",
   768 => x"20286471",
   769 => x"6d292063",
   770 => x"6865636b",
   771 => x"20706173",
   772 => x"7365640a",
   773 => x"00000000",
   774 => x"4c465352",
   775 => x"20636865",
   776 => x"636b2070",
   777 => x"61737365",
   778 => x"642e0a0a",
   779 => x"00000000",
   780 => x"41646472",
   781 => x"65737320",
   782 => x"63686563",
   783 => x"6b207061",
   784 => x"73736564",
   785 => x"2e0a0000",
	others => x"00000000"
);

begin

process (clk)
begin
	if (clk'event and clk = '1') then
		if (from_zpu.memAWriteEnable = '1') and (from_zpu.memBWriteEnable = '1') and (from_zpu.memAAddr=from_zpu.memBAddr) and (from_zpu.memAWrite/=from_zpu.memBWrite) then
			report "write collision" severity failure;
		end if;
	
		if (from_zpu.memAWriteEnable = '1') then
			ram(to_integer(unsigned(from_zpu.memAAddr(maxAddrBitBRAM downto 2)))) := from_zpu.memAWrite;
			to_zpu.memARead <= from_zpu.memAWrite;
		else
			to_zpu.memARead <= ram(to_integer(unsigned(from_zpu.memAAddr(maxAddrBitBRAM downto 2))));
		end if;
	end if;
end process;

process (clk)
begin
	if (clk'event and clk = '1') then
		if (from_zpu.memBWriteEnable = '1') then
			ram(to_integer(unsigned(from_zpu.memBAddr(maxAddrBitBRAM downto 2)))) := from_zpu.memBWrite;
			to_zpu.memBRead <= from_zpu.memBWrite;
		else
			to_zpu.memBRead <= ram(to_integer(unsigned(from_zpu.memBAddr(maxAddrBitBRAM downto 2))));
		end if;
	end if;
end process;


end arch;

