-- ZPU
--
-- Copyright 2004-2008 oharboe - �yvind Harboe - oyvind.harboe@zylin.com
-- Modified by Alastair M. Robinson for the ZPUFlex project.
--
-- The FreeBSD license
-- 
-- Redistribution and use in source and binary forms, with or without
-- modification, are permitted provided that the following conditions
-- are met:
-- 
-- 1. Redistributions of source code must retain the above copyright
--    notice, this list of conditions and the following disclaimer.
-- 2. Redistributions in binary form must reproduce the above
--    copyright notice, this list of conditions and the following
--    disclaimer in the documentation and/or other materials
--    provided with the distribution.
-- 
-- THIS SOFTWARE IS PROVIDED BY THE ZPU PROJECT ``AS IS'' AND ANY
-- EXPRESS OR IMPLIED WARRANTIES, INCLUDING, BUT NOT LIMITED TO,
-- THE IMPLIED WARRANTIES OF MERCHANTABILITY AND FITNESS FOR A
-- PARTICULAR PURPOSE ARE DISCLAIMED. IN NO EVENT SHALL THE
-- ZPU PROJECT OR CONTRIBUTORS BE LIABLE FOR ANY DIRECT,
-- INDIRECT, INCIDENTAL, SPECIAL, EXEMPLARY, OR CONSEQUENTIAL DAMAGES
-- (INCLUDING, BUT NOT LIMITED TO, PROCUREMENT OF SUBSTITUTE GOODS
-- OR SERVICES; LOSS OF USE, DATA, OR PROFITS; OR BUSINESS INTERRUPTION)
-- HOWEVER CAUSED AND ON ANY THEORY OF LIABILITY, WHETHER IN CONTRACT,
-- STRICT LIABILITY, OR TORT (INCLUDING NEGLIGENCE OR OTHERWISE)
-- ARISING IN ANY WAY OUT OF THE USE OF THIS SOFTWARE, EVEN IF
-- ADVISED OF THE POSSIBILITY OF SUCH DAMAGE.
-- 
-- The views and conclusions contained in the software and documentation
-- are those of the authors and should not be interpreted as representing
-- official policies, either expressed or implied, of the ZPU Project.

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;


library work;
use work.zpu_config.all;
use work.zpupkg.all;

entity SDRAMTest_ROM is
generic
	(
		maxAddrBit : integer := maxAddrBitBRAMLimit -- Specify your actual ROM size to save LEs and unnecessary block RAM usage.
	);
port (
	clk : in std_logic;
	areset : in std_logic := '0';
	from_zpu : in ZPU_ToROM;
	to_zpu : out ZPU_FromROM
);
end SDRAMTest_ROM;

architecture arch of SDRAMTest_ROM is

type ram_type is array(natural range 0 to ((2**(maxAddrBit+1))/4)-1) of std_logic_vector(wordSize-1 downto 0);

shared variable ram : ram_type :=
(
     0 => x"0ba08080",
     1 => x"e2040000",
     2 => x"8004a080",
     3 => x"808a0471",
     4 => x"fd060872",
     5 => x"83060981",
     6 => x"05820583",
     7 => x"2b2a83ff",
     8 => x"ff065204",
     9 => x"71fc0608",
    10 => x"72830609",
    11 => x"81058305",
    12 => x"1010102a",
    13 => x"81ff0652",
    14 => x"0471fc06",
    15 => x"080ba080",
    16 => x"8ed47383",
    17 => x"06101005",
    18 => x"08067381",
    19 => x"ff067383",
    20 => x"06098105",
    21 => x"83051010",
    22 => x"102b0772",
    23 => x"fc060c51",
    24 => x"5104a080",
    25 => x"808a0ba0",
    26 => x"808bdc04",
    27 => x"0002c005",
    28 => x"0d0280c4",
    29 => x"05a08095",
    30 => x"c05c5c80",
    31 => x"7c708405",
    32 => x"5e08715f",
    33 => x"5f587d70",
    34 => x"84055f08",
    35 => x"57805a76",
    36 => x"982a7788",
    37 => x"2b585574",
    38 => x"802e8291",
    39 => x"387c802e",
    40 => x"80c23880",
    41 => x"5d7480e4",
    42 => x"2e81b238",
    43 => x"7480e426",
    44 => x"80eb3874",
    45 => x"80e32e80",
    46 => x"c438a551",
    47 => x"a08083b9",
    48 => x"2d7451a0",
    49 => x"8083b92d",
    50 => x"82185881",
    51 => x"1a5a837a",
    52 => x"25ffbc38",
    53 => x"74ffaf38",
    54 => x"7ea08094",
    55 => x"e00c0280",
    56 => x"c0050d04",
    57 => x"74a52e09",
    58 => x"81069a38",
    59 => x"810b811b",
    60 => x"5b5d837a",
    61 => x"25ff9838",
    62 => x"a08081d4",
    63 => x"047b841d",
    64 => x"7108575d",
    65 => x"547451a0",
    66 => x"8083b92d",
    67 => x"8118811b",
    68 => x"5b58837a",
    69 => x"25fef838",
    70 => x"a08081d4",
    71 => x"047480f3",
    72 => x"2e098106",
    73 => x"ff94387b",
    74 => x"841d7108",
    75 => x"70545d5d",
    76 => x"53a08083",
    77 => x"dd2d800b",
    78 => x"ff115452",
    79 => x"807225ff",
    80 => x"8a387a70",
    81 => x"81055c33",
    82 => x"705255a0",
    83 => x"8083b92d",
    84 => x"811873ff",
    85 => x"15555358",
    86 => x"a08082bc",
    87 => x"047b841d",
    88 => x"71087f5c",
    89 => x"555d5287",
    90 => x"56729c2a",
    91 => x"73842b54",
    92 => x"5271802e",
    93 => x"83388159",
    94 => x"b7125471",
    95 => x"89248438",
    96 => x"b0125478",
    97 => x"9438ff16",
    98 => x"56758025",
    99 => x"dc38800b",
   100 => x"ff115452",
   101 => x"a08082bc",
   102 => x"047351a0",
   103 => x"8083b92d",
   104 => x"ff165675",
   105 => x"8025c238",
   106 => x"a080838e",
   107 => x"0477a080",
   108 => x"94e00c02",
   109 => x"80c0050d",
   110 => x"0402f805",
   111 => x"0d7352c0",
   112 => x"0870882a",
   113 => x"70810651",
   114 => x"51517080",
   115 => x"2ef13871",
   116 => x"c00c71a0",
   117 => x"8094e00c",
   118 => x"0288050d",
   119 => x"0402e805",
   120 => x"0d775675",
   121 => x"70840557",
   122 => x"08538054",
   123 => x"72982a73",
   124 => x"882b5452",
   125 => x"71802ea2",
   126 => x"38c00870",
   127 => x"882a7081",
   128 => x"06515151",
   129 => x"70802ef1",
   130 => x"3871c00c",
   131 => x"81158115",
   132 => x"55558374",
   133 => x"25d63871",
   134 => x"ca3874a0",
   135 => x"8094e00c",
   136 => x"0298050d",
   137 => x"0402f405",
   138 => x"0d747652",
   139 => x"53807125",
   140 => x"90387052",
   141 => x"72708405",
   142 => x"5408ff13",
   143 => x"535171f4",
   144 => x"38028c05",
   145 => x"0d0402d4",
   146 => x"050d7c7e",
   147 => x"5c58810b",
   148 => x"a0808ee4",
   149 => x"585a8359",
   150 => x"7608780c",
   151 => x"77087708",
   152 => x"56547375",
   153 => x"2e923877",
   154 => x"08537452",
   155 => x"a0808ef4",
   156 => x"51a08080",
   157 => x"ed2d805a",
   158 => x"7756807b",
   159 => x"2590387a",
   160 => x"55757084",
   161 => x"055708ff",
   162 => x"16565474",
   163 => x"f4387708",
   164 => x"77085656",
   165 => x"75752e92",
   166 => x"38770853",
   167 => x"7452a080",
   168 => x"8fb451a0",
   169 => x"8080ed2d",
   170 => x"805aff19",
   171 => x"84185859",
   172 => x"788025ff",
   173 => x"a33879a0",
   174 => x"8094e00c",
   175 => x"02ac050d",
   176 => x"0402e405",
   177 => x"0d787a55",
   178 => x"56815785",
   179 => x"aad5aad5",
   180 => x"760cfad5",
   181 => x"aad5aa0b",
   182 => x"8c170ccc",
   183 => x"7634b30b",
   184 => x"8f173475",
   185 => x"085372fc",
   186 => x"e2d5aad5",
   187 => x"2e903875",
   188 => x"0852a080",
   189 => x"8ff451a0",
   190 => x"8080ed2d",
   191 => x"80578c16",
   192 => x"085574fa",
   193 => x"d5aad4b3",
   194 => x"2e91388c",
   195 => x"160852a0",
   196 => x"8090b051",
   197 => x"a08080ed",
   198 => x"2d805775",
   199 => x"55807425",
   200 => x"8e387470",
   201 => x"84055608",
   202 => x"ff155553",
   203 => x"73f43875",
   204 => x"085473fc",
   205 => x"e2d5aad5",
   206 => x"2e903875",
   207 => x"0852a080",
   208 => x"90ec51a0",
   209 => x"8080ed2d",
   210 => x"80578c16",
   211 => x"085372fa",
   212 => x"d5aad4b3",
   213 => x"2e91388c",
   214 => x"160852a0",
   215 => x"8091a851",
   216 => x"a08080ed",
   217 => x"2d805776",
   218 => x"a08094e0",
   219 => x"0c029c05",
   220 => x"0d0402c4",
   221 => x"050d605b",
   222 => x"80629080",
   223 => x"8029ff05",
   224 => x"a08091e4",
   225 => x"53405aa0",
   226 => x"8080ed2d",
   227 => x"80e1b357",
   228 => x"80fe5eae",
   229 => x"51a08083",
   230 => x"b92d7610",
   231 => x"70962a81",
   232 => x"06565774",
   233 => x"802e8538",
   234 => x"76810757",
   235 => x"76952a81",
   236 => x"06587780",
   237 => x"2e853876",
   238 => x"81325778",
   239 => x"77077f06",
   240 => x"775e598f",
   241 => x"ffff5876",
   242 => x"bfffff06",
   243 => x"707a3282",
   244 => x"2b7c1151",
   245 => x"57760c76",
   246 => x"1070962a",
   247 => x"81065657",
   248 => x"74802e85",
   249 => x"38768107",
   250 => x"5776952a",
   251 => x"81065574",
   252 => x"802e8538",
   253 => x"76813257",
   254 => x"ff185877",
   255 => x"8025c838",
   256 => x"7c578fff",
   257 => x"ff5876bf",
   258 => x"ffff0670",
   259 => x"7a32822b",
   260 => x"7c057008",
   261 => x"575e5674",
   262 => x"762e80e4",
   263 => x"38807a53",
   264 => x"a08091f4",
   265 => x"525ca080",
   266 => x"80ed2d74",
   267 => x"54755375",
   268 => x"52a08092",
   269 => x"8851a080",
   270 => x"80ed2d7b",
   271 => x"5a761070",
   272 => x"962a8106",
   273 => x"57577580",
   274 => x"2e853876",
   275 => x"81075776",
   276 => x"952a8106",
   277 => x"5574802e",
   278 => x"85387681",
   279 => x"3257ff18",
   280 => x"58778025",
   281 => x"ffa038ff",
   282 => x"1e5e7dfe",
   283 => x"a6388a51",
   284 => x"a08083b9",
   285 => x"2d7ba080",
   286 => x"94e00c02",
   287 => x"bc050d04",
   288 => x"811a5aa0",
   289 => x"8088bd04",
   290 => x"02cc050d",
   291 => x"7e605e58",
   292 => x"815a805b",
   293 => x"80c07a58",
   294 => x"5c85ada9",
   295 => x"89bb780c",
   296 => x"79598156",
   297 => x"97557676",
   298 => x"07822b78",
   299 => x"11515485",
   300 => x"ada989bb",
   301 => x"740c7510",
   302 => x"ff165656",
   303 => x"748025e6",
   304 => x"38761081",
   305 => x"1a5a5798",
   306 => x"7925d738",
   307 => x"7756807d",
   308 => x"2590387c",
   309 => x"55757084",
   310 => x"055708ff",
   311 => x"16565474",
   312 => x"f4388157",
   313 => x"ff8787a5",
   314 => x"c3780c97",
   315 => x"5976822b",
   316 => x"78117008",
   317 => x"5f56567c",
   318 => x"ff8787a5",
   319 => x"c32e80c7",
   320 => x"38740854",
   321 => x"7385ada9",
   322 => x"89bb2e92",
   323 => x"38807508",
   324 => x"547653a0",
   325 => x"8092b052",
   326 => x"5aa08080",
   327 => x"ed2d7610",
   328 => x"ff1a5a57",
   329 => x"788025c5",
   330 => x"387a822b",
   331 => x"5675ad38",
   332 => x"7b52a080",
   333 => x"92d051a0",
   334 => x"8080ed2d",
   335 => x"7ba08094",
   336 => x"e00c02b4",
   337 => x"050d047a",
   338 => x"77077710",
   339 => x"ff1b5b58",
   340 => x"5b788025",
   341 => x"ff9738a0",
   342 => x"808aa904",
   343 => x"7552a080",
   344 => x"938c51a0",
   345 => x"8080ed2d",
   346 => x"75992a81",
   347 => x"32810670",
   348 => x"09810571",
   349 => x"07700970",
   350 => x"9f2c7d06",
   351 => x"79109fff",
   352 => x"fffc0660",
   353 => x"812a415a",
   354 => x"5d575859",
   355 => x"75da3879",
   356 => x"09810570",
   357 => x"7b079f2a",
   358 => x"55567bbf",
   359 => x"26843873",
   360 => x"9a388170",
   361 => x"53a08092",
   362 => x"d0525ca0",
   363 => x"8080ed2d",
   364 => x"7ba08094",
   365 => x"e00c02b4",
   366 => x"050d04a0",
   367 => x"8093a451",
   368 => x"a08080ed",
   369 => x"2d7b52a0",
   370 => x"8092d051",
   371 => x"a08080ed",
   372 => x"2d7ba080",
   373 => x"94e00c02",
   374 => x"b4050d04",
   375 => x"02dc050d",
   376 => x"810ba080",
   377 => x"8ee45858",
   378 => x"83597608",
   379 => x"800c8008",
   380 => x"77085654",
   381 => x"73752e92",
   382 => x"38800853",
   383 => x"7452a080",
   384 => x"8ef451a0",
   385 => x"8080ed2d",
   386 => x"80588070",
   387 => x"57557570",
   388 => x"84055708",
   389 => x"81165654",
   390 => x"a0807524",
   391 => x"f1388008",
   392 => x"77085656",
   393 => x"75752e92",
   394 => x"38800853",
   395 => x"7452a080",
   396 => x"8fb451a0",
   397 => x"8080ed2d",
   398 => x"8058ff19",
   399 => x"84185859",
   400 => x"788025ff",
   401 => x"a5387780",
   402 => x"2e8b38a0",
   403 => x"8093f051",
   404 => x"a08080ed",
   405 => x"2d815785",
   406 => x"aad5aad5",
   407 => x"0b800cfa",
   408 => x"d5aad5aa",
   409 => x"0b8c0ccc",
   410 => x"0b8034b3",
   411 => x"0b8f3480",
   412 => x"085574fc",
   413 => x"e2d5aad5",
   414 => x"2e903880",
   415 => x"0852a080",
   416 => x"8ff451a0",
   417 => x"8080ed2d",
   418 => x"80578c08",
   419 => x"5877fad5",
   420 => x"aad4b32e",
   421 => x"90388c08",
   422 => x"52a08090",
   423 => x"b051a080",
   424 => x"80ed2d80",
   425 => x"57807057",
   426 => x"55757084",
   427 => x"05570881",
   428 => x"165654a0",
   429 => x"807524f1",
   430 => x"38800859",
   431 => x"78fce2d5",
   432 => x"aad52e90",
   433 => x"38800852",
   434 => x"a08090ec",
   435 => x"51a08080",
   436 => x"ed2d8057",
   437 => x"8c085473",
   438 => x"fad5aad4",
   439 => x"b32e80dd",
   440 => x"388c0852",
   441 => x"a08091a8",
   442 => x"51a08080",
   443 => x"ed2da080",
   444 => x"528051a0",
   445 => x"8089882d",
   446 => x"a08094e0",
   447 => x"0854a080",
   448 => x"94e00880",
   449 => x"2e8b38a0",
   450 => x"80949451",
   451 => x"a08080ed",
   452 => x"2d735280",
   453 => x"51a08086",
   454 => x"f22da080",
   455 => x"94e00880",
   456 => x"2efdbd38",
   457 => x"a08094ac",
   458 => x"51a08080",
   459 => x"ed2d810b",
   460 => x"a0808ee4",
   461 => x"58588359",
   462 => x"a0808bea",
   463 => x"0476802e",
   464 => x"ffac38a0",
   465 => x"8094c451",
   466 => x"a08080ed",
   467 => x"2da0808d",
   468 => x"ee040000",
   469 => x"00ffffff",
   470 => x"ff00ffff",
   471 => x"ffff00ff",
   472 => x"ffffff00",
   473 => x"00000000",
   474 => x"55555555",
   475 => x"aaaaaaaa",
   476 => x"ffffffff",
   477 => x"53616e69",
   478 => x"74792063",
   479 => x"6865636b",
   480 => x"20666169",
   481 => x"6c656420",
   482 => x"28626566",
   483 => x"6f726520",
   484 => x"63616368",
   485 => x"65207265",
   486 => x"66726573",
   487 => x"6829206f",
   488 => x"6e203078",
   489 => x"25642028",
   490 => x"676f7420",
   491 => x"30782564",
   492 => x"290a0000",
   493 => x"53616e69",
   494 => x"74792063",
   495 => x"6865636b",
   496 => x"20666169",
   497 => x"6c656420",
   498 => x"28616674",
   499 => x"65722063",
   500 => x"61636865",
   501 => x"20726566",
   502 => x"72657368",
   503 => x"29206f6e",
   504 => x"20307825",
   505 => x"64202867",
   506 => x"6f742030",
   507 => x"78256429",
   508 => x"0a000000",
   509 => x"42797465",
   510 => x"20636865",
   511 => x"636b2066",
   512 => x"61696c65",
   513 => x"64202862",
   514 => x"65666f72",
   515 => x"65206361",
   516 => x"63686520",
   517 => x"72656672",
   518 => x"65736829",
   519 => x"20617420",
   520 => x"30202867",
   521 => x"6f742030",
   522 => x"78256429",
   523 => x"0a000000",
   524 => x"42797465",
   525 => x"20636865",
   526 => x"636b2066",
   527 => x"61696c65",
   528 => x"64202862",
   529 => x"65666f72",
   530 => x"65206361",
   531 => x"63686520",
   532 => x"72656672",
   533 => x"65736829",
   534 => x"20617420",
   535 => x"33202867",
   536 => x"6f742030",
   537 => x"78256429",
   538 => x"0a000000",
   539 => x"42797465",
   540 => x"20636865",
   541 => x"636b2066",
   542 => x"61696c65",
   543 => x"64202861",
   544 => x"66746572",
   545 => x"20636163",
   546 => x"68652072",
   547 => x"65667265",
   548 => x"73682920",
   549 => x"61742030",
   550 => x"2028676f",
   551 => x"74203078",
   552 => x"2564290a",
   553 => x"00000000",
   554 => x"42797465",
   555 => x"20636865",
   556 => x"636b2066",
   557 => x"61696c65",
   558 => x"64202861",
   559 => x"66746572",
   560 => x"20636163",
   561 => x"68652072",
   562 => x"65667265",
   563 => x"73682920",
   564 => x"61742033",
   565 => x"2028676f",
   566 => x"74203078",
   567 => x"2564290a",
   568 => x"00000000",
   569 => x"43686563",
   570 => x"6b696e67",
   571 => x"206d656d",
   572 => x"6f727900",
   573 => x"30782564",
   574 => x"20676f6f",
   575 => x"64207265",
   576 => x"6164732c",
   577 => x"20000000",
   578 => x"4572726f",
   579 => x"72206174",
   580 => x"20307825",
   581 => x"642c2065",
   582 => x"78706563",
   583 => x"74656420",
   584 => x"30782564",
   585 => x"2c20676f",
   586 => x"74203078",
   587 => x"25640a00",
   588 => x"42616420",
   589 => x"64617461",
   590 => x"20666f75",
   591 => x"6e642061",
   592 => x"74203078",
   593 => x"25642028",
   594 => x"30782564",
   595 => x"290a0000",
   596 => x"53445241",
   597 => x"4d207369",
   598 => x"7a652028",
   599 => x"61737375",
   600 => x"6d696e67",
   601 => x"206e6f20",
   602 => x"61646472",
   603 => x"65737320",
   604 => x"6661756c",
   605 => x"74732920",
   606 => x"69732030",
   607 => x"78256420",
   608 => x"6d656761",
   609 => x"62797465",
   610 => x"730a0000",
   611 => x"416c6961",
   612 => x"73657320",
   613 => x"666f756e",
   614 => x"64206174",
   615 => x"20307825",
   616 => x"640a0000",
   617 => x"28416c69",
   618 => x"61736573",
   619 => x"2070726f",
   620 => x"6261626c",
   621 => x"79207369",
   622 => x"6d706c79",
   623 => x"20696e64",
   624 => x"69636174",
   625 => x"65207468",
   626 => x"61742052",
   627 => x"414d0a69",
   628 => x"7320736d",
   629 => x"616c6c65",
   630 => x"72207468",
   631 => x"616e2036",
   632 => x"34206d65",
   633 => x"67616279",
   634 => x"74657329",
   635 => x"0a000000",
   636 => x"46697273",
   637 => x"74207374",
   638 => x"61676520",
   639 => x"73616e69",
   640 => x"74792063",
   641 => x"6865636b",
   642 => x"20706173",
   643 => x"7365642e",
   644 => x"0a000000",
   645 => x"41646472",
   646 => x"65737320",
   647 => x"63686563",
   648 => x"6b207061",
   649 => x"73736564",
   650 => x"2e0a0000",
   651 => x"4c465352",
   652 => x"20636865",
   653 => x"636b2070",
   654 => x"61737365",
   655 => x"642e0a0a",
   656 => x"00000000",
   657 => x"42797465",
   658 => x"20286471",
   659 => x"6d292063",
   660 => x"6865636b",
   661 => x"20706173",
   662 => x"7365640a",
   663 => x"00000000",
	others => x"00000000"
);

begin

process (clk)
begin
	if (clk'event and clk = '1') then
		if (from_zpu.memAWriteEnable = '1') and (from_zpu.memBWriteEnable = '1') and (from_zpu.memAAddr=from_zpu.memBAddr) and (from_zpu.memAWrite/=from_zpu.memBWrite) then
			report "write collision" severity failure;
		end if;
	
		if (from_zpu.memAWriteEnable = '1') then
			ram(to_integer(unsigned(from_zpu.memAAddr(maxAddrBit downto 2)))) := from_zpu.memAWrite;
			to_zpu.memARead <= from_zpu.memAWrite;
		else
			to_zpu.memARead <= ram(to_integer(unsigned(from_zpu.memAAddr(maxAddrBit downto 2))));
		end if;
	end if;
end process;

process (clk)
begin
	if (clk'event and clk = '1') then
		if (from_zpu.memBWriteEnable = '1') then
			ram(to_integer(unsigned(from_zpu.memBAddr(maxAddrBit downto 2)))) := from_zpu.memBWrite;
			to_zpu.memBRead <= from_zpu.memBWrite;
		else
			to_zpu.memBRead <= ram(to_integer(unsigned(from_zpu.memBAddr(maxAddrBit downto 2))));
		end if;
	end if;
end process;


end arch;

