-- ZPU
--
-- Copyright 2004-2008 oharboe - �yvind Harboe - oyvind.harboe@zylin.com
-- Modified by Alastair M. Robinson for the ZPUFlex project.
--
-- The FreeBSD license
-- 
-- Redistribution and use in source and binary forms, with or without
-- modification, are permitted provided that the following conditions
-- are met:
-- 
-- 1. Redistributions of source code must retain the above copyright
--    notice, this list of conditions and the following disclaimer.
-- 2. Redistributions in binary form must reproduce the above
--    copyright notice, this list of conditions and the following
--    disclaimer in the documentation and/or other materials
--    provided with the distribution.
-- 
-- THIS SOFTWARE IS PROVIDED BY THE ZPU PROJECT ``AS IS'' AND ANY
-- EXPRESS OR IMPLIED WARRANTIES, INCLUDING, BUT NOT LIMITED TO,
-- THE IMPLIED WARRANTIES OF MERCHANTABILITY AND FITNESS FOR A
-- PARTICULAR PURPOSE ARE DISCLAIMED. IN NO EVENT SHALL THE
-- ZPU PROJECT OR CONTRIBUTORS BE LIABLE FOR ANY DIRECT,
-- INDIRECT, INCIDENTAL, SPECIAL, EXEMPLARY, OR CONSEQUENTIAL DAMAGES
-- (INCLUDING, BUT NOT LIMITED TO, PROCUREMENT OF SUBSTITUTE GOODS
-- OR SERVICES; LOSS OF USE, DATA, OR PROFITS; OR BUSINESS INTERRUPTION)
-- HOWEVER CAUSED AND ON ANY THEORY OF LIABILITY, WHETHER IN CONTRACT,
-- STRICT LIABILITY, OR TORT (INCLUDING NEGLIGENCE OR OTHERWISE)
-- ARISING IN ANY WAY OUT OF THE USE OF THIS SOFTWARE, EVEN IF
-- ADVISED OF THE POSSIBILITY OF SUCH DAMAGE.
-- 
-- The views and conclusions contained in the software and documentation
-- are those of the authors and should not be interpreted as representing
-- official policies, either expressed or implied, of the ZPU Project.

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;


library work;
use work.zpu_config.all;
use work.zpupkg.all;

entity Interrupt_ROM is
generic
	(
		maxAddrBit : integer := maxAddrBitBRAMLimit -- Specify your actual ROM size to save LEs and unnecessary block RAM usage.
	);
port (
	clk : in std_logic;
	areset : in std_logic := '0';
	from_zpu : in ZPU_ToROM;
	to_zpu : out ZPU_FromROM
);
end Interrupt_ROM;

architecture arch of Interrupt_ROM is

type ram_type is array(natural range 0 to ((2**(maxAddrBit+1))/4)-1) of std_logic_vector(wordSize-1 downto 0);

shared variable ram : ram_type :=
(
     0 => x"0b0b0b88",
     1 => x"dd040000",
     2 => x"00000000",
     3 => x"00000000",
     4 => x"00000000",
     5 => x"00000000",
     6 => x"00000000",
     7 => x"00000000",
     8 => x"88088c08",
     9 => x"90080b0b",
    10 => x"0b88e708",
    11 => x"2d900c8c",
    12 => x"0c880c04",
    13 => x"00000000",
    14 => x"00000000",
    15 => x"00000000",
    16 => x"71fd0608",
    17 => x"72830609",
    18 => x"81058205",
    19 => x"832b2a83",
    20 => x"ffff0652",
    21 => x"04000000",
    22 => x"00000000",
    23 => x"00000000",
    24 => x"71fd0608",
    25 => x"83ffff73",
    26 => x"83060981",
    27 => x"05820583",
    28 => x"2b2b0906",
    29 => x"7383ffff",
    30 => x"0b0b0b0b",
    31 => x"83a50400",
    32 => x"72098105",
    33 => x"72057373",
    34 => x"09060906",
    35 => x"73097306",
    36 => x"070a8106",
    37 => x"53510400",
    38 => x"00000000",
    39 => x"00000000",
    40 => x"72722473",
    41 => x"732e0753",
    42 => x"51040000",
    43 => x"00000000",
    44 => x"00000000",
    45 => x"00000000",
    46 => x"00000000",
    47 => x"00000000",
    48 => x"71737109",
    49 => x"71068106",
    50 => x"09810572",
    51 => x"0a100a72",
    52 => x"0a100a31",
    53 => x"050a8106",
    54 => x"51515351",
    55 => x"04000000",
    56 => x"72722673",
    57 => x"732e0753",
    58 => x"51040000",
    59 => x"00000000",
    60 => x"00000000",
    61 => x"00000000",
    62 => x"00000000",
    63 => x"00000000",
    64 => x"00000000",
    65 => x"00000000",
    66 => x"00000000",
    67 => x"00000000",
    68 => x"00000000",
    69 => x"00000000",
    70 => x"00000000",
    71 => x"00000000",
    72 => x"0b0b0b88",
    73 => x"ba040000",
    74 => x"00000000",
    75 => x"00000000",
    76 => x"00000000",
    77 => x"00000000",
    78 => x"00000000",
    79 => x"00000000",
    80 => x"720a722b",
    81 => x"0a535104",
    82 => x"00000000",
    83 => x"00000000",
    84 => x"00000000",
    85 => x"00000000",
    86 => x"00000000",
    87 => x"00000000",
    88 => x"72729f06",
    89 => x"0981050b",
    90 => x"0b0b889f",
    91 => x"05040000",
    92 => x"00000000",
    93 => x"00000000",
    94 => x"00000000",
    95 => x"00000000",
    96 => x"72722aff",
    97 => x"739f062a",
    98 => x"0974090a",
    99 => x"8106ff05",
   100 => x"06075351",
   101 => x"04000000",
   102 => x"00000000",
   103 => x"00000000",
   104 => x"71715351",
   105 => x"04067383",
   106 => x"06098105",
   107 => x"8205832b",
   108 => x"0b2b0772",
   109 => x"fc060c51",
   110 => x"51040000",
   111 => x"00000000",
   112 => x"72098105",
   113 => x"72050970",
   114 => x"81050906",
   115 => x"0a810653",
   116 => x"51040000",
   117 => x"00000000",
   118 => x"00000000",
   119 => x"00000000",
   120 => x"72098105",
   121 => x"72050970",
   122 => x"81050906",
   123 => x"0a098106",
   124 => x"53510400",
   125 => x"00000000",
   126 => x"00000000",
   127 => x"00000000",
   128 => x"71098105",
   129 => x"52040000",
   130 => x"00000000",
   131 => x"00000000",
   132 => x"00000000",
   133 => x"00000000",
   134 => x"00000000",
   135 => x"00000000",
   136 => x"72720981",
   137 => x"05055351",
   138 => x"04000000",
   139 => x"00000000",
   140 => x"00000000",
   141 => x"00000000",
   142 => x"00000000",
   143 => x"00000000",
   144 => x"72097206",
   145 => x"73730906",
   146 => x"07535104",
   147 => x"00000000",
   148 => x"00000000",
   149 => x"00000000",
   150 => x"00000000",
   151 => x"00000000",
   152 => x"71fc0608",
   153 => x"72830609",
   154 => x"81058305",
   155 => x"1010102a",
   156 => x"81ff0652",
   157 => x"04000000",
   158 => x"00000000",
   159 => x"00000000",
   160 => x"71fc0608",
   161 => x"0b0b0b91",
   162 => x"98738306",
   163 => x"10100508",
   164 => x"060b0b0b",
   165 => x"88a20400",
   166 => x"00000000",
   167 => x"00000000",
   168 => x"88088c08",
   169 => x"90087575",
   170 => x"0b0b0b8d",
   171 => x"9c2d5050",
   172 => x"88085690",
   173 => x"0c8c0c88",
   174 => x"0c510400",
   175 => x"00000000",
   176 => x"88088c08",
   177 => x"90087575",
   178 => x"0b0b0b8e",
   179 => x"ce2d5050",
   180 => x"88085690",
   181 => x"0c8c0c88",
   182 => x"0c510400",
   183 => x"00000000",
   184 => x"72097081",
   185 => x"0509060a",
   186 => x"8106ff05",
   187 => x"70547106",
   188 => x"73097274",
   189 => x"05ff0506",
   190 => x"07515151",
   191 => x"04000000",
   192 => x"72097081",
   193 => x"0509060a",
   194 => x"098106ff",
   195 => x"05705471",
   196 => x"06730972",
   197 => x"7405ff05",
   198 => x"06075151",
   199 => x"51040000",
   200 => x"05ff0504",
   201 => x"00000000",
   202 => x"00000000",
   203 => x"00000000",
   204 => x"00000000",
   205 => x"00000000",
   206 => x"00000000",
   207 => x"00000000",
   208 => x"04000000",
   209 => x"00000000",
   210 => x"00000000",
   211 => x"00000000",
   212 => x"00000000",
   213 => x"00000000",
   214 => x"00000000",
   215 => x"00000000",
   216 => x"71810552",
   217 => x"04000000",
   218 => x"00000000",
   219 => x"00000000",
   220 => x"00000000",
   221 => x"00000000",
   222 => x"00000000",
   223 => x"00000000",
   224 => x"00000000",
   225 => x"00000000",
   226 => x"00000000",
   227 => x"00000000",
   228 => x"00000000",
   229 => x"00000000",
   230 => x"00000000",
   231 => x"00000000",
   232 => x"02840572",
   233 => x"10100552",
   234 => x"04000000",
   235 => x"00000000",
   236 => x"00000000",
   237 => x"00000000",
   238 => x"00000000",
   239 => x"00000000",
   240 => x"00000000",
   241 => x"00000000",
   242 => x"00000000",
   243 => x"00000000",
   244 => x"00000000",
   245 => x"00000000",
   246 => x"00000000",
   247 => x"00000000",
   248 => x"717105ff",
   249 => x"05715351",
   250 => x"020d0400",
   251 => x"00000000",
   252 => x"00000000",
   253 => x"00000000",
   254 => x"00000000",
   255 => x"00000000",
   256 => x"10101010",
   257 => x"10101010",
   258 => x"10101010",
   259 => x"10101010",
   260 => x"10101010",
   261 => x"10101010",
   262 => x"10101010",
   263 => x"10101053",
   264 => x"51047381",
   265 => x"ff067383",
   266 => x"06098105",
   267 => x"83051010",
   268 => x"102b0772",
   269 => x"fc060c51",
   270 => x"51047272",
   271 => x"80728106",
   272 => x"ff050972",
   273 => x"06057110",
   274 => x"52720a10",
   275 => x"0a5372ed",
   276 => x"38515153",
   277 => x"51040000",
   278 => x"800488da",
   279 => x"0488da0b",
   280 => x"8cb90404",
   281 => x"00000000",
   282 => x"000463f1",
   283 => x"3d0d923d",
   284 => x"0b0b0b92",
   285 => x"bc5c5680",
   286 => x"76708405",
   287 => x"5808715f",
   288 => x"5f577d70",
   289 => x"84055f08",
   290 => x"5a805c79",
   291 => x"982a7a88",
   292 => x"2b5b5574",
   293 => x"8638765f",
   294 => x"81f8397c",
   295 => x"802e81d2",
   296 => x"38805d74",
   297 => x"80e42e9b",
   298 => x"387480e4",
   299 => x"268b3874",
   300 => x"80e32e81",
   301 => x"8a388191",
   302 => x"397480f3",
   303 => x"2e80ef38",
   304 => x"81873975",
   305 => x"84177108",
   306 => x"0b0b0b92",
   307 => x"bc0b0b0b",
   308 => x"0b91ec61",
   309 => x"5d585c52",
   310 => x"5753728e",
   311 => x"38b00b0b",
   312 => x"0b0b91ec",
   313 => x"34811454",
   314 => x"ae398a52",
   315 => x"72518387",
   316 => x"3f88080b",
   317 => x"0b0b91a8",
   318 => x"05337470",
   319 => x"81055634",
   320 => x"8a527251",
   321 => x"82cc3f88",
   322 => x"08538808",
   323 => x"dd38730b",
   324 => x"0b0b91ec",
   325 => x"2e9138ff",
   326 => x"14547333",
   327 => x"79708105",
   328 => x"5b348118",
   329 => x"58e83980",
   330 => x"79347754",
   331 => x"ab397584",
   332 => x"17710870",
   333 => x"545d5753",
   334 => x"80fe3f7c",
   335 => x"549a3975",
   336 => x"84177108",
   337 => x"575753b6",
   338 => x"39a55180",
   339 => x"cc3f7451",
   340 => x"80c73f82",
   341 => x"1757ae39",
   342 => x"73ff1555",
   343 => x"53807325",
   344 => x"a4387a70",
   345 => x"81055c33",
   346 => x"705255ad",
   347 => x"3f811757",
   348 => x"e73974a5",
   349 => x"2e098106",
   350 => x"8538815d",
   351 => x"88397451",
   352 => x"983f8117",
   353 => x"57811c5c",
   354 => x"837c25fd",
   355 => x"fe3874fd",
   356 => x"f1387e88",
   357 => x"0c913d0d",
   358 => x"04ff3d0d",
   359 => x"7352c008",
   360 => x"70882a70",
   361 => x"81065151",
   362 => x"5170802e",
   363 => x"f13871c0",
   364 => x"0c71880c",
   365 => x"833d0d04",
   366 => x"fb3d0d77",
   367 => x"55747084",
   368 => x"05560853",
   369 => x"80547298",
   370 => x"2a73882b",
   371 => x"54527180",
   372 => x"2ea238c0",
   373 => x"0870882a",
   374 => x"70810651",
   375 => x"51517080",
   376 => x"2ef13871",
   377 => x"c00c8116",
   378 => x"81155556",
   379 => x"837425d6",
   380 => x"3871ca38",
   381 => x"75880c87",
   382 => x"3d0d0471",
   383 => x"88e70c04",
   384 => x"ffb00888",
   385 => x"0c04810b",
   386 => x"ffb00c04",
   387 => x"800bffb0",
   388 => x"0c04ff3d",
   389 => x"0df63fe8",
   390 => x"3f92fc08",
   391 => x"81327092",
   392 => x"fc0c5271",
   393 => x"802e8638",
   394 => x"91bc5184",
   395 => x"3991c851",
   396 => x"ff863fd2",
   397 => x"3f833d0d",
   398 => x"04803d0d",
   399 => x"800b92fc",
   400 => x"0c91d451",
   401 => x"fef23f8c",
   402 => x"9251ffaf",
   403 => x"3fffb73f",
   404 => x"ff399408",
   405 => x"02940cfd",
   406 => x"3d0d8053",
   407 => x"94088c05",
   408 => x"08529408",
   409 => x"88050851",
   410 => x"82de3f88",
   411 => x"0870880c",
   412 => x"54853d0d",
   413 => x"940c0494",
   414 => x"0802940c",
   415 => x"fd3d0d81",
   416 => x"5394088c",
   417 => x"05085294",
   418 => x"08880508",
   419 => x"5182b93f",
   420 => x"88087088",
   421 => x"0c54853d",
   422 => x"0d940c04",
   423 => x"94080294",
   424 => x"0cf93d0d",
   425 => x"800b9408",
   426 => x"fc050c94",
   427 => x"08880508",
   428 => x"8025ab38",
   429 => x"94088805",
   430 => x"08309408",
   431 => x"88050c80",
   432 => x"0b9408f4",
   433 => x"050c9408",
   434 => x"fc050888",
   435 => x"38810b94",
   436 => x"08f4050c",
   437 => x"9408f405",
   438 => x"089408fc",
   439 => x"050c9408",
   440 => x"8c050880",
   441 => x"25ab3894",
   442 => x"088c0508",
   443 => x"3094088c",
   444 => x"050c800b",
   445 => x"9408f005",
   446 => x"0c9408fc",
   447 => x"05088838",
   448 => x"810b9408",
   449 => x"f0050c94",
   450 => x"08f00508",
   451 => x"9408fc05",
   452 => x"0c805394",
   453 => x"088c0508",
   454 => x"52940888",
   455 => x"05085181",
   456 => x"a73f8808",
   457 => x"709408f8",
   458 => x"050c5494",
   459 => x"08fc0508",
   460 => x"802e8c38",
   461 => x"9408f805",
   462 => x"08309408",
   463 => x"f8050c94",
   464 => x"08f80508",
   465 => x"70880c54",
   466 => x"893d0d94",
   467 => x"0c049408",
   468 => x"02940cfb",
   469 => x"3d0d800b",
   470 => x"9408fc05",
   471 => x"0c940888",
   472 => x"05088025",
   473 => x"93389408",
   474 => x"88050830",
   475 => x"94088805",
   476 => x"0c810b94",
   477 => x"08fc050c",
   478 => x"94088c05",
   479 => x"0880258c",
   480 => x"3894088c",
   481 => x"05083094",
   482 => x"088c050c",
   483 => x"81539408",
   484 => x"8c050852",
   485 => x"94088805",
   486 => x"0851ad3f",
   487 => x"88087094",
   488 => x"08f8050c",
   489 => x"549408fc",
   490 => x"0508802e",
   491 => x"8c389408",
   492 => x"f8050830",
   493 => x"9408f805",
   494 => x"0c9408f8",
   495 => x"05087088",
   496 => x"0c54873d",
   497 => x"0d940c04",
   498 => x"94080294",
   499 => x"0cfd3d0d",
   500 => x"810b9408",
   501 => x"fc050c80",
   502 => x"0b9408f8",
   503 => x"050c9408",
   504 => x"8c050894",
   505 => x"08880508",
   506 => x"27ac3894",
   507 => x"08fc0508",
   508 => x"802ea338",
   509 => x"800b9408",
   510 => x"8c050824",
   511 => x"99389408",
   512 => x"8c050810",
   513 => x"94088c05",
   514 => x"0c9408fc",
   515 => x"05081094",
   516 => x"08fc050c",
   517 => x"c9399408",
   518 => x"fc050880",
   519 => x"2e80c938",
   520 => x"94088c05",
   521 => x"08940888",
   522 => x"050826a1",
   523 => x"38940888",
   524 => x"05089408",
   525 => x"8c050831",
   526 => x"94088805",
   527 => x"0c9408f8",
   528 => x"05089408",
   529 => x"fc050807",
   530 => x"9408f805",
   531 => x"0c9408fc",
   532 => x"0508812a",
   533 => x"9408fc05",
   534 => x"0c94088c",
   535 => x"0508812a",
   536 => x"94088c05",
   537 => x"0cffaf39",
   538 => x"94089005",
   539 => x"08802e8f",
   540 => x"38940888",
   541 => x"05087094",
   542 => x"08f4050c",
   543 => x"518d3994",
   544 => x"08f80508",
   545 => x"709408f4",
   546 => x"050c5194",
   547 => x"08f40508",
   548 => x"880c853d",
   549 => x"0d940c04",
   550 => x"00ffffff",
   551 => x"ff00ffff",
   552 => x"ffff00ff",
   553 => x"ffffff00",
   554 => x"30313233",
   555 => x"34353637",
   556 => x"38394142",
   557 => x"43444546",
   558 => x"00000000",
   559 => x"5469636b",
   560 => x"2e2e2e0a",
   561 => x"00000000",
   562 => x"546f636b",
   563 => x"2e2e2e0a",
   564 => x"00000000",
   565 => x"456e6162",
   566 => x"6c696e67",
   567 => x"20696e74",
   568 => x"65727275",
   569 => x"7074732e",
   570 => x"2e2e0a00",
	others => x"00000000"
);

begin

process (clk)
begin
	if (clk'event and clk = '1') then
		if (from_zpu.memAWriteEnable = '1') and (from_zpu.memBWriteEnable = '1') and (from_zpu.memAAddr=from_zpu.memBAddr) and (from_zpu.memAWrite/=from_zpu.memBWrite) then
			report "write collision" severity failure;
		end if;
	
		if (from_zpu.memAWriteEnable = '1') then
			ram(to_integer(unsigned(from_zpu.memAAddr(maxAddrBit downto 2)))) := from_zpu.memAWrite;
			to_zpu.memARead <= from_zpu.memAWrite;
		else
			to_zpu.memARead <= ram(to_integer(unsigned(from_zpu.memAAddr(maxAddrBit downto 2))));
		end if;
	end if;
end process;

process (clk)
begin
	if (clk'event and clk = '1') then
		if (from_zpu.memBWriteEnable = '1') then
			ram(to_integer(unsigned(from_zpu.memBAddr(maxAddrBit downto 2)))) := from_zpu.memBWrite;
			to_zpu.memBRead <= from_zpu.memBWrite;
		else
			to_zpu.memBRead <= ram(to_integer(unsigned(from_zpu.memBAddr(maxAddrBit downto 2))));
		end if;
	end if;
end process;


end arch;

