-- ZPU
--
-- Copyright 2004-2008 oharboe - �yvind Harboe - oyvind.harboe@zylin.com
-- Modified by Alastair M. Robinson for the ZPUFlex project.
--
-- The FreeBSD license
-- 
-- Redistribution and use in source and binary forms, with or without
-- modification, are permitted provided that the following conditions
-- are met:
-- 
-- 1. Redistributions of source code must retain the above copyright
--    notice, this list of conditions and the following disclaimer.
-- 2. Redistributions in binary form must reproduce the above
--    copyright notice, this list of conditions and the following
--    disclaimer in the documentation and/or other materials
--    provided with the distribution.
-- 
-- THIS SOFTWARE IS PROVIDED BY THE ZPU PROJECT ``AS IS'' AND ANY
-- EXPRESS OR IMPLIED WARRANTIES, INCLUDING, BUT NOT LIMITED TO,
-- THE IMPLIED WARRANTIES OF MERCHANTABILITY AND FITNESS FOR A
-- PARTICULAR PURPOSE ARE DISCLAIMED. IN NO EVENT SHALL THE
-- ZPU PROJECT OR CONTRIBUTORS BE LIABLE FOR ANY DIRECT,
-- INDIRECT, INCIDENTAL, SPECIAL, EXEMPLARY, OR CONSEQUENTIAL DAMAGES
-- (INCLUDING, BUT NOT LIMITED TO, PROCUREMENT OF SUBSTITUTE GOODS
-- OR SERVICES; LOSS OF USE, DATA, OR PROFITS; OR BUSINESS INTERRUPTION)
-- HOWEVER CAUSED AND ON ANY THEORY OF LIABILITY, WHETHER IN CONTRACT,
-- STRICT LIABILITY, OR TORT (INCLUDING NEGLIGENCE OR OTHERWISE)
-- ARISING IN ANY WAY OUT OF THE USE OF THIS SOFTWARE, EVEN IF
-- ADVISED OF THE POSSIBILITY OF SUCH DAMAGE.
-- 
-- The views and conclusions contained in the software and documentation
-- are those of the authors and should not be interpreted as representing
-- official policies, either expressed or implied, of the ZPU Project.

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;


library work;
use work.zpu_config.all;
use work.zpupkg.all;

entity VGATest_ROM is
generic
	(
		maxAddrBitBRAM : integer := maxAddrBitBRAMLimit -- Specify your actual ROM size to save LEs and unnecessary block RAM usage.
	);
port (
	clk : in std_logic;
	areset : in std_logic := '0';
	from_zpu : in ZPU_ToROM;
	to_zpu : out ZPU_FromROM
);
end VGATest_ROM;

architecture arch of VGATest_ROM is

type ram_type is array(natural range 0 to ((2**(maxAddrBitBRAM+1))/4)-1) of std_logic_vector(wordSize-1 downto 0);

shared variable ram : ram_type :=
(
     0 => x"84808080",
     1 => x"ed040000",
     2 => x"00000000",
     3 => x"84808080",
     4 => x"880d8004",
     5 => x"84808080",
     6 => x"940471fd",
     7 => x"06087283",
     8 => x"06098105",
     9 => x"8205832b",
    10 => x"2a83ffff",
    11 => x"06520471",
    12 => x"fc060872",
    13 => x"83060981",
    14 => x"05830510",
    15 => x"10102a81",
    16 => x"ff065204",
    17 => x"71fc0608",
    18 => x"84808091",
    19 => x"d0738306",
    20 => x"10100508",
    21 => x"067381ff",
    22 => x"06738306",
    23 => x"09810583",
    24 => x"05101010",
    25 => x"2b0772fc",
    26 => x"060c5151",
    27 => x"04028405",
    28 => x"84808080",
    29 => x"880c8480",
    30 => x"8080940b",
    31 => x"84808085",
    32 => x"86040000",
    33 => x"02c0050d",
    34 => x"0280c405",
    35 => x"84808098",
    36 => x"bc5c5c80",
    37 => x"7c708405",
    38 => x"5e08715f",
    39 => x"5f587d70",
    40 => x"84055f08",
    41 => x"57805976",
    42 => x"982a7788",
    43 => x"2b585574",
    44 => x"802e82ae",
    45 => x"387c802e",
    46 => x"80c53880",
    47 => x"5d7480e4",
    48 => x"2e81c038",
    49 => x"7480e426",
    50 => x"80f13874",
    51 => x"80e32e80",
    52 => x"c838a551",
    53 => x"84808084",
    54 => x"962d7451",
    55 => x"84808084",
    56 => x"962d8218",
    57 => x"58811959",
    58 => x"837925ff",
    59 => x"ba3874ff",
    60 => x"ad387e84",
    61 => x"808097dc",
    62 => x"0c0280c0",
    63 => x"050d0474",
    64 => x"a52e0981",
    65 => x"069b3881",
    66 => x"0b811a5a",
    67 => x"5d837925",
    68 => x"ff953884",
    69 => x"808081ee",
    70 => x"047b841d",
    71 => x"7108575d",
    72 => x"54745184",
    73 => x"80808496",
    74 => x"2d811881",
    75 => x"1a5a5883",
    76 => x"7925fef3",
    77 => x"38848080",
    78 => x"81ee0474",
    79 => x"80f32e09",
    80 => x"8106ff8e",
    81 => x"387b841d",
    82 => x"71087054",
    83 => x"5d5d5384",
    84 => x"808084bb",
    85 => x"2d800bff",
    86 => x"11545280",
    87 => x"7225ff85",
    88 => x"387a7081",
    89 => x"055c8480",
    90 => x"8080af2d",
    91 => x"70525584",
    92 => x"80808496",
    93 => x"2d811873",
    94 => x"ff155553",
    95 => x"58848080",
    96 => x"82db047b",
    97 => x"841d7108",
    98 => x"7f5d555d",
    99 => x"52807324",
   100 => x"80f13872",
   101 => x"802e80d7",
   102 => x"38875672",
   103 => x"9c2a7384",
   104 => x"2b545271",
   105 => x"802e8338",
   106 => x"815ab712",
   107 => x"54718924",
   108 => x"8438b012",
   109 => x"54799538",
   110 => x"ff165675",
   111 => x"8025dc38",
   112 => x"800bff11",
   113 => x"54528480",
   114 => x"8082db04",
   115 => x"73518480",
   116 => x"8084962d",
   117 => x"ff165675",
   118 => x"8025c038",
   119 => x"84808083",
   120 => x"c0047784",
   121 => x"808097dc",
   122 => x"0c0280c0",
   123 => x"050d04b0",
   124 => x"51848080",
   125 => x"84962d80",
   126 => x"0bff1154",
   127 => x"52848080",
   128 => x"82db04ad",
   129 => x"51848080",
   130 => x"84962d72",
   131 => x"09810553",
   132 => x"84808083",
   133 => x"930402f8",
   134 => x"050d7352",
   135 => x"c0087088",
   136 => x"2a708106",
   137 => x"51515170",
   138 => x"802ef138",
   139 => x"71c00c71",
   140 => x"84808097",
   141 => x"dc0c0288",
   142 => x"050d0402",
   143 => x"e8050d80",
   144 => x"78575575",
   145 => x"70840557",
   146 => x"08538054",
   147 => x"72982a73",
   148 => x"882b5452",
   149 => x"71802ea2",
   150 => x"38c00870",
   151 => x"882a7081",
   152 => x"06515151",
   153 => x"70802ef1",
   154 => x"3871c00c",
   155 => x"81158115",
   156 => x"55558374",
   157 => x"25d63871",
   158 => x"ca387484",
   159 => x"808097dc",
   160 => x"0c029805",
   161 => x"0d0402dc",
   162 => x"050d8052",
   163 => x"8480800b",
   164 => x"fc800c81",
   165 => x"12705559",
   166 => x"84808056",
   167 => x"805584fe",
   168 => x"53811483",
   169 => x"ffff0670",
   170 => x"77708405",
   171 => x"590cfe14",
   172 => x"54547280",
   173 => x"25eb3881",
   174 => x"155583df",
   175 => x"7525df38",
   176 => x"80578055",
   177 => x"84fe53fc",
   178 => x"8008fe14",
   179 => x"54527280",
   180 => x"25f53881",
   181 => x"155583df",
   182 => x"7525e938",
   183 => x"811757b1",
   184 => x"7725df38",
   185 => x"80587555",
   186 => x"805784fe",
   187 => x"53811483",
   188 => x"ffff0670",
   189 => x"76708405",
   190 => x"580cfe14",
   191 => x"54547280",
   192 => x"25eb3881",
   193 => x"175783df",
   194 => x"7725df38",
   195 => x"81185893",
   196 => x"7825d338",
   197 => x"81195280",
   198 => x"51848080",
   199 => x"8e8f2d84",
   200 => x"80808593",
   201 => x"0402f405",
   202 => x"0d747652",
   203 => x"53807125",
   204 => x"90387052",
   205 => x"72708405",
   206 => x"5408ff13",
   207 => x"535171f4",
   208 => x"38028c05",
   209 => x"0d0402d4",
   210 => x"050d7c7e",
   211 => x"5c58810b",
   212 => x"84808091",
   213 => x"e0585a83",
   214 => x"59760878",
   215 => x"0c770877",
   216 => x"08565473",
   217 => x"752e9438",
   218 => x"77085374",
   219 => x"52848080",
   220 => x"91f05184",
   221 => x"80808184",
   222 => x"2d805a77",
   223 => x"56807b25",
   224 => x"90387a55",
   225 => x"75708405",
   226 => x"5708ff16",
   227 => x"565474f4",
   228 => x"38770877",
   229 => x"08565675",
   230 => x"752e9438",
   231 => x"77085374",
   232 => x"52848080",
   233 => x"92b05184",
   234 => x"80808184",
   235 => x"2d805aff",
   236 => x"19841858",
   237 => x"59788025",
   238 => x"ff9f3879",
   239 => x"84808097",
   240 => x"dc0c02ac",
   241 => x"050d0402",
   242 => x"e4050d78",
   243 => x"7a555681",
   244 => x"5785aad5",
   245 => x"aad5760c",
   246 => x"fad5aad5",
   247 => x"aa0b8c17",
   248 => x"0ccc7684",
   249 => x"808080c4",
   250 => x"2db30b8f",
   251 => x"17848080",
   252 => x"80c42d75",
   253 => x"085372fc",
   254 => x"e2d5aad5",
   255 => x"2e923875",
   256 => x"08528480",
   257 => x"8092f051",
   258 => x"84808081",
   259 => x"842d8057",
   260 => x"8c160855",
   261 => x"74fad5aa",
   262 => x"d4b32e93",
   263 => x"388c1608",
   264 => x"52848080",
   265 => x"93ac5184",
   266 => x"80808184",
   267 => x"2d805775",
   268 => x"55807425",
   269 => x"8e387470",
   270 => x"84055608",
   271 => x"ff155553",
   272 => x"73f43875",
   273 => x"085473fc",
   274 => x"e2d5aad5",
   275 => x"2e923875",
   276 => x"08528480",
   277 => x"8093e851",
   278 => x"84808081",
   279 => x"842d8057",
   280 => x"8c160853",
   281 => x"72fad5aa",
   282 => x"d4b32e93",
   283 => x"388c1608",
   284 => x"52848080",
   285 => x"94a45184",
   286 => x"80808184",
   287 => x"2d805776",
   288 => x"84808097",
   289 => x"dc0c029c",
   290 => x"050d0402",
   291 => x"c4050d60",
   292 => x"5b806290",
   293 => x"808029ff",
   294 => x"05848080",
   295 => x"94e05340",
   296 => x"5a848080",
   297 => x"81842d80",
   298 => x"e1b35780",
   299 => x"fe5eae51",
   300 => x"84808084",
   301 => x"962d7610",
   302 => x"70962a81",
   303 => x"06565774",
   304 => x"802e8538",
   305 => x"76810757",
   306 => x"76952a81",
   307 => x"06587780",
   308 => x"2e853876",
   309 => x"81325778",
   310 => x"77077f06",
   311 => x"775e598f",
   312 => x"ffff5876",
   313 => x"bfffff06",
   314 => x"707a3282",
   315 => x"2b7c1151",
   316 => x"57760c76",
   317 => x"1070962a",
   318 => x"81065657",
   319 => x"74802e85",
   320 => x"38768107",
   321 => x"5776952a",
   322 => x"81065574",
   323 => x"802e8538",
   324 => x"76813257",
   325 => x"ff185877",
   326 => x"8025c838",
   327 => x"7c578fff",
   328 => x"ff5876bf",
   329 => x"ffff0670",
   330 => x"7a32822b",
   331 => x"7c057008",
   332 => x"575e5674",
   333 => x"762e80ea",
   334 => x"38807a53",
   335 => x"84808094",
   336 => x"f0525c84",
   337 => x"80808184",
   338 => x"2d745475",
   339 => x"53755284",
   340 => x"80809584",
   341 => x"51848080",
   342 => x"81842d7b",
   343 => x"5a761070",
   344 => x"962a8106",
   345 => x"57577580",
   346 => x"2e853876",
   347 => x"81075776",
   348 => x"952a8106",
   349 => x"5574802e",
   350 => x"85387681",
   351 => x"3257ff18",
   352 => x"58778025",
   353 => x"ff9c38ff",
   354 => x"1e5e7dfe",
   355 => x"a1388a51",
   356 => x"84808084",
   357 => x"962d7b84",
   358 => x"808097dc",
   359 => x"0c02bc05",
   360 => x"0d04811a",
   361 => x"5a848080",
   362 => x"8add0402",
   363 => x"cc050d7e",
   364 => x"605e5881",
   365 => x"5a805b80",
   366 => x"c07a585c",
   367 => x"85ada989",
   368 => x"bb780c79",
   369 => x"59815697",
   370 => x"55767607",
   371 => x"822b7811",
   372 => x"515485ad",
   373 => x"a989bb74",
   374 => x"0c7510ff",
   375 => x"16565674",
   376 => x"8025e638",
   377 => x"7610811a",
   378 => x"5a579879",
   379 => x"25d73877",
   380 => x"56807d25",
   381 => x"90387c55",
   382 => x"75708405",
   383 => x"5708ff16",
   384 => x"565474f4",
   385 => x"388157ff",
   386 => x"8787a5c3",
   387 => x"780c9759",
   388 => x"76822b78",
   389 => x"1170085f",
   390 => x"56567cff",
   391 => x"8787a5c3",
   392 => x"2e80cc38",
   393 => x"74085473",
   394 => x"85ada989",
   395 => x"bb2e9438",
   396 => x"80750854",
   397 => x"76538480",
   398 => x"8095ac52",
   399 => x"5a848080",
   400 => x"81842d76",
   401 => x"10ff1a5a",
   402 => x"57788025",
   403 => x"c3387a82",
   404 => x"2b5675b1",
   405 => x"387b5284",
   406 => x"808095cc",
   407 => x"51848080",
   408 => x"81842d7b",
   409 => x"84808097",
   410 => x"dc0c02b4",
   411 => x"050d047a",
   412 => x"77077710",
   413 => x"ff1b5b58",
   414 => x"5b788025",
   415 => x"ff923884",
   416 => x"80808cce",
   417 => x"04755284",
   418 => x"80809688",
   419 => x"51848080",
   420 => x"81842d75",
   421 => x"992a8132",
   422 => x"81067009",
   423 => x"81057107",
   424 => x"7009709f",
   425 => x"2c7d0679",
   426 => x"109fffff",
   427 => x"fc066081",
   428 => x"2a415a5d",
   429 => x"57585975",
   430 => x"da387909",
   431 => x"8105707b",
   432 => x"079f2a55",
   433 => x"567bbf26",
   434 => x"8438739d",
   435 => x"38817053",
   436 => x"84808095",
   437 => x"cc525c84",
   438 => x"80808184",
   439 => x"2d7b8480",
   440 => x"8097dc0c",
   441 => x"02b4050d",
   442 => x"04848080",
   443 => x"96a05184",
   444 => x"80808184",
   445 => x"2d7b5284",
   446 => x"808095cc",
   447 => x"51848080",
   448 => x"81842d7b",
   449 => x"84808097",
   450 => x"dc0c02b4",
   451 => x"050d0402",
   452 => x"d4050d7c",
   453 => x"57817084",
   454 => x"808091e0",
   455 => x"5b595b83",
   456 => x"5a780877",
   457 => x"0c760879",
   458 => x"08565473",
   459 => x"752e9438",
   460 => x"76085374",
   461 => x"52848080",
   462 => x"91f05184",
   463 => x"80808184",
   464 => x"2d805876",
   465 => x"569fff55",
   466 => x"75708405",
   467 => x"5708ff16",
   468 => x"56547480",
   469 => x"25f23876",
   470 => x"08790856",
   471 => x"5675752e",
   472 => x"94387608",
   473 => x"53745284",
   474 => x"808092b0",
   475 => x"51848080",
   476 => x"81842d80",
   477 => x"58ff1a84",
   478 => x"1a5a5a79",
   479 => x"8025ffa1",
   480 => x"387781fd",
   481 => x"38775b81",
   482 => x"5885aad5",
   483 => x"aad5770c",
   484 => x"fad5aad5",
   485 => x"aa0b8c18",
   486 => x"0ccc7784",
   487 => x"808080c4",
   488 => x"2db30b8f",
   489 => x"18848080",
   490 => x"80c42d76",
   491 => x"085574fc",
   492 => x"e2d5aad5",
   493 => x"2e923876",
   494 => x"08528480",
   495 => x"8092f051",
   496 => x"84808081",
   497 => x"842d8058",
   498 => x"8c170859",
   499 => x"78fad5aa",
   500 => x"d4b32e93",
   501 => x"388c1708",
   502 => x"52848080",
   503 => x"93ac5184",
   504 => x"80808184",
   505 => x"2d805876",
   506 => x"569fff55",
   507 => x"75708405",
   508 => x"5708ff16",
   509 => x"56547480",
   510 => x"25f23876",
   511 => x"085a79fc",
   512 => x"e2d5aad5",
   513 => x"2e923876",
   514 => x"08528480",
   515 => x"8093e851",
   516 => x"84808081",
   517 => x"842d8058",
   518 => x"8c170854",
   519 => x"73fad5aa",
   520 => x"d4b32e80",
   521 => x"ee388c17",
   522 => x"08528480",
   523 => x"8094a451",
   524 => x"84808081",
   525 => x"842d8058",
   526 => x"775ba080",
   527 => x"52765184",
   528 => x"80808bab",
   529 => x"2d848080",
   530 => x"97dc0854",
   531 => x"84808097",
   532 => x"dc0880e9",
   533 => x"38848080",
   534 => x"97dc085b",
   535 => x"73527651",
   536 => x"84808089",
   537 => x"8b2d8480",
   538 => x"8097dc08",
   539 => x"be388480",
   540 => x"8097dc08",
   541 => x"5b7a8480",
   542 => x"8097dc0c",
   543 => x"02ac050d",
   544 => x"04848080",
   545 => x"96ec5184",
   546 => x"80808184",
   547 => x"2d848080",
   548 => x"8f870477",
   549 => x"802effa0",
   550 => x"38848080",
   551 => x"97905184",
   552 => x"80808184",
   553 => x"2d848080",
   554 => x"90ba0484",
   555 => x"808097ac",
   556 => x"51848080",
   557 => x"81842d84",
   558 => x"808090f5",
   559 => x"04848080",
   560 => x"97c45184",
   561 => x"80808184",
   562 => x"2d848080",
   563 => x"90dc0400",
   564 => x"00ffffff",
   565 => x"ff00ffff",
   566 => x"ffff00ff",
   567 => x"ffffff00",
   568 => x"00000000",
   569 => x"55555555",
   570 => x"aaaaaaaa",
   571 => x"ffffffff",
   572 => x"53616e69",
   573 => x"74792063",
   574 => x"6865636b",
   575 => x"20666169",
   576 => x"6c656420",
   577 => x"28626566",
   578 => x"6f726520",
   579 => x"63616368",
   580 => x"65207265",
   581 => x"66726573",
   582 => x"6829206f",
   583 => x"6e203078",
   584 => x"25642028",
   585 => x"676f7420",
   586 => x"30782564",
   587 => x"290a0000",
   588 => x"53616e69",
   589 => x"74792063",
   590 => x"6865636b",
   591 => x"20666169",
   592 => x"6c656420",
   593 => x"28616674",
   594 => x"65722063",
   595 => x"61636865",
   596 => x"20726566",
   597 => x"72657368",
   598 => x"29206f6e",
   599 => x"20307825",
   600 => x"64202867",
   601 => x"6f742030",
   602 => x"78256429",
   603 => x"0a000000",
   604 => x"42797465",
   605 => x"20636865",
   606 => x"636b2066",
   607 => x"61696c65",
   608 => x"64202862",
   609 => x"65666f72",
   610 => x"65206361",
   611 => x"63686520",
   612 => x"72656672",
   613 => x"65736829",
   614 => x"20617420",
   615 => x"30202867",
   616 => x"6f742030",
   617 => x"78256429",
   618 => x"0a000000",
   619 => x"42797465",
   620 => x"20636865",
   621 => x"636b2066",
   622 => x"61696c65",
   623 => x"64202862",
   624 => x"65666f72",
   625 => x"65206361",
   626 => x"63686520",
   627 => x"72656672",
   628 => x"65736829",
   629 => x"20617420",
   630 => x"33202867",
   631 => x"6f742030",
   632 => x"78256429",
   633 => x"0a000000",
   634 => x"42797465",
   635 => x"20636865",
   636 => x"636b2066",
   637 => x"61696c65",
   638 => x"64202861",
   639 => x"66746572",
   640 => x"20636163",
   641 => x"68652072",
   642 => x"65667265",
   643 => x"73682920",
   644 => x"61742030",
   645 => x"2028676f",
   646 => x"74203078",
   647 => x"2564290a",
   648 => x"00000000",
   649 => x"42797465",
   650 => x"20636865",
   651 => x"636b2066",
   652 => x"61696c65",
   653 => x"64202861",
   654 => x"66746572",
   655 => x"20636163",
   656 => x"68652072",
   657 => x"65667265",
   658 => x"73682920",
   659 => x"61742033",
   660 => x"2028676f",
   661 => x"74203078",
   662 => x"2564290a",
   663 => x"00000000",
   664 => x"43686563",
   665 => x"6b696e67",
   666 => x"206d656d",
   667 => x"6f727900",
   668 => x"30782564",
   669 => x"20676f6f",
   670 => x"64207265",
   671 => x"6164732c",
   672 => x"20000000",
   673 => x"4572726f",
   674 => x"72206174",
   675 => x"20307825",
   676 => x"642c2065",
   677 => x"78706563",
   678 => x"74656420",
   679 => x"30782564",
   680 => x"2c20676f",
   681 => x"74203078",
   682 => x"25640a00",
   683 => x"42616420",
   684 => x"64617461",
   685 => x"20666f75",
   686 => x"6e642061",
   687 => x"74203078",
   688 => x"25642028",
   689 => x"30782564",
   690 => x"290a0000",
   691 => x"53445241",
   692 => x"4d207369",
   693 => x"7a652028",
   694 => x"61737375",
   695 => x"6d696e67",
   696 => x"206e6f20",
   697 => x"61646472",
   698 => x"65737320",
   699 => x"6661756c",
   700 => x"74732920",
   701 => x"69732030",
   702 => x"78256420",
   703 => x"6d656761",
   704 => x"62797465",
   705 => x"730a0000",
   706 => x"416c6961",
   707 => x"73657320",
   708 => x"666f756e",
   709 => x"64206174",
   710 => x"20307825",
   711 => x"640a0000",
   712 => x"28416c69",
   713 => x"61736573",
   714 => x"2070726f",
   715 => x"6261626c",
   716 => x"79207369",
   717 => x"6d706c79",
   718 => x"20696e64",
   719 => x"69636174",
   720 => x"65207468",
   721 => x"61742052",
   722 => x"414d0a69",
   723 => x"7320736d",
   724 => x"616c6c65",
   725 => x"72207468",
   726 => x"616e2036",
   727 => x"34206d65",
   728 => x"67616279",
   729 => x"74657329",
   730 => x"0a000000",
   731 => x"46697273",
   732 => x"74207374",
   733 => x"61676520",
   734 => x"73616e69",
   735 => x"74792063",
   736 => x"6865636b",
   737 => x"20706173",
   738 => x"7365642e",
   739 => x"0a000000",
   740 => x"42797465",
   741 => x"20286471",
   742 => x"6d292063",
   743 => x"6865636b",
   744 => x"20706173",
   745 => x"7365640a",
   746 => x"00000000",
   747 => x"4c465352",
   748 => x"20636865",
   749 => x"636b2070",
   750 => x"61737365",
   751 => x"642e0a0a",
   752 => x"00000000",
   753 => x"41646472",
   754 => x"65737320",
   755 => x"63686563",
   756 => x"6b207061",
   757 => x"73736564",
   758 => x"2e0a0000",
	others => x"00000000"
);

begin

process (clk)
begin
	if (clk'event and clk = '1') then
		if (from_zpu.memAWriteEnable = '1') and (from_zpu.memBWriteEnable = '1') and (from_zpu.memAAddr=from_zpu.memBAddr) and (from_zpu.memAWrite/=from_zpu.memBWrite) then
			report "write collision" severity failure;
		end if;
	
		if (from_zpu.memAWriteEnable = '1') then
			ram(to_integer(unsigned(from_zpu.memAAddr(maxAddrBitBRAM downto 2)))) := from_zpu.memAWrite;
			to_zpu.memARead <= from_zpu.memAWrite;
		else
			to_zpu.memARead <= ram(to_integer(unsigned(from_zpu.memAAddr(maxAddrBitBRAM downto 2))));
		end if;
	end if;
end process;

process (clk)
begin
	if (clk'event and clk = '1') then
		if (from_zpu.memBWriteEnable = '1') then
			ram(to_integer(unsigned(from_zpu.memBAddr(maxAddrBitBRAM downto 2)))) := from_zpu.memBWrite;
			to_zpu.memBRead <= from_zpu.memBWrite;
		else
			to_zpu.memBRead <= ram(to_integer(unsigned(from_zpu.memBAddr(maxAddrBitBRAM downto 2))));
		end if;
	end if;
end process;


end arch;

