-- ZPU
--
-- Copyright 2004-2008 oharboe - �yvind Harboe - oyvind.harboe@zylin.com
-- Modified by Alastair M. Robinson for the ZPUFlex project.
--
-- The FreeBSD license
-- 
-- Redistribution and use in source and binary forms, with or without
-- modification, are permitted provided that the following conditions
-- are met:
-- 
-- 1. Redistributions of source code must retain the above copyright
--    notice, this list of conditions and the following disclaimer.
-- 2. Redistributions in binary form must reproduce the above
--    copyright notice, this list of conditions and the following
--    disclaimer in the documentation and/or other materials
--    provided with the distribution.
-- 
-- THIS SOFTWARE IS PROVIDED BY THE ZPU PROJECT ``AS IS'' AND ANY
-- EXPRESS OR IMPLIED WARRANTIES, INCLUDING, BUT NOT LIMITED TO,
-- THE IMPLIED WARRANTIES OF MERCHANTABILITY AND FITNESS FOR A
-- PARTICULAR PURPOSE ARE DISCLAIMED. IN NO EVENT SHALL THE
-- ZPU PROJECT OR CONTRIBUTORS BE LIABLE FOR ANY DIRECT,
-- INDIRECT, INCIDENTAL, SPECIAL, EXEMPLARY, OR CONSEQUENTIAL DAMAGES
-- (INCLUDING, BUT NOT LIMITED TO, PROCUREMENT OF SUBSTITUTE GOODS
-- OR SERVICES; LOSS OF USE, DATA, OR PROFITS; OR BUSINESS INTERRUPTION)
-- HOWEVER CAUSED AND ON ANY THEORY OF LIABILITY, WHETHER IN CONTRACT,
-- STRICT LIABILITY, OR TORT (INCLUDING NEGLIGENCE OR OTHERWISE)
-- ARISING IN ANY WAY OUT OF THE USE OF THIS SOFTWARE, EVEN IF
-- ADVISED OF THE POSSIBILITY OF SUCH DAMAGE.
-- 
-- The views and conclusions contained in the software and documentation
-- are those of the authors and should not be interpreted as representing
-- official policies, either expressed or implied, of the ZPU Project.

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;


library work;
use work.zpu_config.all;
use work.zpupkg.all;

entity SDBootstrap_ROM is
generic
	(
		maxAddrBitBRAM : integer := maxAddrBitBRAMLimit -- Specify your actual ROM size to save LEs and unnecessary block RAM usage.
	);
port (
	clk : in std_logic;
	areset : in std_logic := '0';
	from_zpu : in ZPU_ToROM;
	to_zpu : out ZPU_FromROM
);
end SDBootstrap_ROM;

architecture arch of SDBootstrap_ROM is

type ram_type is array(natural range 0 to ((2**(maxAddrBitBRAM+1))/4)-1) of std_logic_vector(wordSize-1 downto 0);

shared variable ram : ram_type :=
(
     0 => x"0ba08080",
     1 => x"ec040000",
     2 => x"00000000",
     3 => x"0ba08080",
     4 => x"880d8004",
     5 => x"a0808094",
     6 => x"0471fd06",
     7 => x"08728306",
     8 => x"09810582",
     9 => x"05832b2a",
    10 => x"83ffff06",
    11 => x"520471fc",
    12 => x"06087283",
    13 => x"06098105",
    14 => x"83051010",
    15 => x"102a81ff",
    16 => x"06520471",
    17 => x"fc06080b",
    18 => x"a0809e88",
    19 => x"73830610",
    20 => x"10050806",
    21 => x"7381ff06",
    22 => x"73830609",
    23 => x"81058305",
    24 => x"1010102b",
    25 => x"0772fc06",
    26 => x"0c515104",
    27 => x"0284050b",
    28 => x"a0808088",
    29 => x"0ca08080",
    30 => x"940ba080",
    31 => x"8cba0400",
    32 => x"0002c405",
    33 => x"0d0280c0",
    34 => x"0583ffe0",
    35 => x"e05b5680",
    36 => x"76708405",
    37 => x"5808715e",
    38 => x"5e577c70",
    39 => x"84055e08",
    40 => x"58805b77",
    41 => x"982a7888",
    42 => x"2b595372",
    43 => x"8838765e",
    44 => x"a08083aa",
    45 => x"047b802e",
    46 => x"81ca3880",
    47 => x"5c7280e4",
    48 => x"2e9f3872",
    49 => x"80e4268d",
    50 => x"387280e3",
    51 => x"2e80ee38",
    52 => x"a08082ca",
    53 => x"047280f3",
    54 => x"2e80cc38",
    55 => x"a08082ca",
    56 => x"04758417",
    57 => x"71087e5c",
    58 => x"56575287",
    59 => x"55739c2a",
    60 => x"74842b55",
    61 => x"5271802e",
    62 => x"83388159",
    63 => x"89722589",
    64 => x"38b71252",
    65 => x"a080828c",
    66 => x"04b01252",
    67 => x"78802e88",
    68 => x"387151a0",
    69 => x"8083b52d",
    70 => x"ff155574",
    71 => x"8025ce38",
    72 => x"8054a080",
    73 => x"82e00475",
    74 => x"84177108",
    75 => x"70545c57",
    76 => x"52a08083",
    77 => x"d92d7b54",
    78 => x"a08082e0",
    79 => x"04758417",
    80 => x"71085557",
    81 => x"52a08083",
    82 => x"9304a551",
    83 => x"a08083b5",
    84 => x"2d7251a0",
    85 => x"8083b52d",
    86 => x"821757a0",
    87 => x"80839d04",
    88 => x"73ff1555",
    89 => x"52807225",
    90 => x"b4387970",
    91 => x"81055ba0",
    92 => x"8080ae2d",
    93 => x"705253a0",
    94 => x"8083b52d",
    95 => x"811757a0",
    96 => x"8082e004",
    97 => x"72a52e09",
    98 => x"81068838",
    99 => x"815ca080",
   100 => x"839d0472",
   101 => x"51a08083",
   102 => x"b52d8117",
   103 => x"57811b5b",
   104 => x"837b25fd",
   105 => x"fe3872fd",
   106 => x"f1387d83",
   107 => x"ffe0800c",
   108 => x"02bc050d",
   109 => x"0402f805",
   110 => x"0d7352c0",
   111 => x"0870882a",
   112 => x"70810651",
   113 => x"51517080",
   114 => x"2ef13871",
   115 => x"c00c7183",
   116 => x"ffe0800c",
   117 => x"0288050d",
   118 => x"0402e805",
   119 => x"0d807857",
   120 => x"55757084",
   121 => x"05570853",
   122 => x"80547298",
   123 => x"2a73882b",
   124 => x"54527180",
   125 => x"2ea238c0",
   126 => x"0870882a",
   127 => x"70810651",
   128 => x"51517080",
   129 => x"2ef13871",
   130 => x"c00c8115",
   131 => x"81155555",
   132 => x"837425d6",
   133 => x"3871ca38",
   134 => x"7483ffe0",
   135 => x"800c0298",
   136 => x"050d0402",
   137 => x"f4050d74",
   138 => x"767181ff",
   139 => x"06d40c53",
   140 => x"5383fff1",
   141 => x"a0088538",
   142 => x"71892b52",
   143 => x"71982ad4",
   144 => x"0c71902a",
   145 => x"7081ff06",
   146 => x"d40c5171",
   147 => x"882a7081",
   148 => x"ff06d40c",
   149 => x"517181ff",
   150 => x"06d40c72",
   151 => x"902a7081",
   152 => x"ff06d40c",
   153 => x"51d40870",
   154 => x"81ff0651",
   155 => x"5182b8bf",
   156 => x"527081ff",
   157 => x"2e098106",
   158 => x"943881ff",
   159 => x"0bd40cd4",
   160 => x"087081ff",
   161 => x"06ff1454",
   162 => x"515171e5",
   163 => x"387083ff",
   164 => x"e0800c02",
   165 => x"8c050d04",
   166 => x"02fc050d",
   167 => x"81c75181",
   168 => x"ff0bd40c",
   169 => x"ff115170",
   170 => x"8025f438",
   171 => x"0284050d",
   172 => x"0402f005",
   173 => x"0da08085",
   174 => x"982d819c",
   175 => x"9f538052",
   176 => x"87fc80f7",
   177 => x"51a08084",
   178 => x"a32d83ff",
   179 => x"e0800854",
   180 => x"83ffe080",
   181 => x"08812e09",
   182 => x"8106ab38",
   183 => x"81ff0bd4",
   184 => x"0c820a52",
   185 => x"849c80e9",
   186 => x"51a08084",
   187 => x"a32d83ff",
   188 => x"e080088d",
   189 => x"3881ff0b",
   190 => x"d40c7353",
   191 => x"a080868d",
   192 => x"04a08085",
   193 => x"982dff13",
   194 => x"5372ffb2",
   195 => x"387283ff",
   196 => x"e0800c02",
   197 => x"90050d04",
   198 => x"02f4050d",
   199 => x"81ff0bd4",
   200 => x"0ca0809e",
   201 => x"9851a080",
   202 => x"83d92d93",
   203 => x"53805287",
   204 => x"fc80c151",
   205 => x"a08084a3",
   206 => x"2d83ffe0",
   207 => x"80088d38",
   208 => x"81ff0bd4",
   209 => x"0c8153a0",
   210 => x"8086d704",
   211 => x"a0808598",
   212 => x"2dff1353",
   213 => x"72d73872",
   214 => x"83ffe080",
   215 => x"0c028c05",
   216 => x"0d0402f0",
   217 => x"050da080",
   218 => x"85982d83",
   219 => x"aa52849c",
   220 => x"80c851a0",
   221 => x"8084a32d",
   222 => x"83ffe080",
   223 => x"0883ffe0",
   224 => x"800853a0",
   225 => x"809ea452",
   226 => x"54a08081",
   227 => x"812d7381",
   228 => x"2e098106",
   229 => x"9038d808",
   230 => x"7083ffff",
   231 => x"06545472",
   232 => x"83aa2ea3",
   233 => x"38a08086",
   234 => x"982da080",
   235 => x"87c00481",
   236 => x"54a08088",
   237 => x"eb04a080",
   238 => x"9ebc51a0",
   239 => x"8081812d",
   240 => x"8054a080",
   241 => x"88eb0473",
   242 => x"52a0809e",
   243 => x"d851a080",
   244 => x"81812d81",
   245 => x"ff0bd40c",
   246 => x"b153a080",
   247 => x"85b12d83",
   248 => x"ffe08008",
   249 => x"802e80f4",
   250 => x"38805287",
   251 => x"fc80fa51",
   252 => x"a08084a3",
   253 => x"2d83ffe0",
   254 => x"800880d0",
   255 => x"3883ffe0",
   256 => x"800852a0",
   257 => x"809ef051",
   258 => x"a0808181",
   259 => x"2d81ff0b",
   260 => x"d40cd408",
   261 => x"81ff0670",
   262 => x"53a0809e",
   263 => x"fc5254a0",
   264 => x"8081812d",
   265 => x"81ff0bd4",
   266 => x"0c81ff0b",
   267 => x"d40c81ff",
   268 => x"0bd40c81",
   269 => x"ff0bd40c",
   270 => x"73862a70",
   271 => x"81067056",
   272 => x"51537280",
   273 => x"2ea538a0",
   274 => x"8087af04",
   275 => x"83ffe080",
   276 => x"0852a080",
   277 => x"9ef051a0",
   278 => x"8081812d",
   279 => x"72822efe",
   280 => x"d538ff13",
   281 => x"5372fef2",
   282 => x"38725473",
   283 => x"83ffe080",
   284 => x"0c029005",
   285 => x"0d0402f4",
   286 => x"050d810b",
   287 => x"83fff1a0",
   288 => x"0cd00870",
   289 => x"8f2a7081",
   290 => x"06515153",
   291 => x"72f33872",
   292 => x"d00ca080",
   293 => x"85982dd0",
   294 => x"08708f2a",
   295 => x"70810651",
   296 => x"515372f3",
   297 => x"38810bd0",
   298 => x"0c875380",
   299 => x"5284d480",
   300 => x"c051a080",
   301 => x"84a32d83",
   302 => x"ffe08008",
   303 => x"812e9638",
   304 => x"72822e09",
   305 => x"81068838",
   306 => x"8053a080",
   307 => x"8a8d04ff",
   308 => x"135372d7",
   309 => x"38a08086",
   310 => x"e22d83ff",
   311 => x"e0800883",
   312 => x"fff1a00c",
   313 => x"815287fc",
   314 => x"80d051a0",
   315 => x"8084a32d",
   316 => x"81ff0bd4",
   317 => x"0cd00870",
   318 => x"8f2a7081",
   319 => x"06515153",
   320 => x"72f33872",
   321 => x"d00c81ff",
   322 => x"0bd40c81",
   323 => x"537283ff",
   324 => x"e0800c02",
   325 => x"8c050d04",
   326 => x"800b83ff",
   327 => x"e0800c04",
   328 => x"02e0050d",
   329 => x"797b5757",
   330 => x"805881ff",
   331 => x"0bd40cd0",
   332 => x"08708f2a",
   333 => x"70810651",
   334 => x"515473f3",
   335 => x"3882810b",
   336 => x"d00c81ff",
   337 => x"0bd40c76",
   338 => x"5287fc80",
   339 => x"d151a080",
   340 => x"84a32d80",
   341 => x"dbc6df55",
   342 => x"83ffe080",
   343 => x"08802e98",
   344 => x"3883ffe0",
   345 => x"80085376",
   346 => x"52a0809f",
   347 => x"8c51a080",
   348 => x"81812da0",
   349 => x"808bc404",
   350 => x"81ff0bd4",
   351 => x"0cd40870",
   352 => x"81ff0651",
   353 => x"547381fe",
   354 => x"2e098106",
   355 => x"9b3880ff",
   356 => x"55d80876",
   357 => x"70840558",
   358 => x"0cff1555",
   359 => x"748025f1",
   360 => x"388158a0",
   361 => x"808bae04",
   362 => x"ff155574",
   363 => x"cb3881ff",
   364 => x"0bd40cd0",
   365 => x"08708f2a",
   366 => x"70810651",
   367 => x"515473f3",
   368 => x"3873d00c",
   369 => x"7783ffe0",
   370 => x"800c02a0",
   371 => x"050d0402",
   372 => x"f4050d74",
   373 => x"70882a83",
   374 => x"fe800670",
   375 => x"72982a07",
   376 => x"72882b87",
   377 => x"fc808006",
   378 => x"73982b81",
   379 => x"f00a0671",
   380 => x"73070783",
   381 => x"ffe0800c",
   382 => x"56515351",
   383 => x"028c050d",
   384 => x"0402f805",
   385 => x"0d028e05",
   386 => x"a08080ae",
   387 => x"2d74982b",
   388 => x"71902b07",
   389 => x"70902c83",
   390 => x"ffe0800c",
   391 => x"52520288",
   392 => x"050d0402",
   393 => x"f8050d73",
   394 => x"70902b71",
   395 => x"902a0783",
   396 => x"ffe0800c",
   397 => x"52028805",
   398 => x"0d0402ec",
   399 => x"050d800b",
   400 => x"fc800ca0",
   401 => x"809fac51",
   402 => x"a08083d9",
   403 => x"2da08088",
   404 => x"f62d83ff",
   405 => x"e0800880",
   406 => x"2e81e638",
   407 => x"a0809fc4",
   408 => x"51a08083",
   409 => x"d92da080",
   410 => x"8f9f2d83",
   411 => x"ffe1a052",
   412 => x"a0809fdc",
   413 => x"51a0809b",
   414 => x"a82d83ff",
   415 => x"e0800880",
   416 => x"2e81be38",
   417 => x"83ffe1a0",
   418 => x"0ba0809f",
   419 => x"e85254a0",
   420 => x"8083d92d",
   421 => x"80557370",
   422 => x"810555a0",
   423 => x"8080ae2d",
   424 => x"5372a02e",
   425 => x"80de3872",
   426 => x"a32e80fd",
   427 => x"387280c7",
   428 => x"2e098106",
   429 => x"8b38a080",
   430 => x"808c2da0",
   431 => x"808de004",
   432 => x"728a2e09",
   433 => x"81068b38",
   434 => x"a0808094",
   435 => x"2da0808d",
   436 => x"e0047280",
   437 => x"cc2e0981",
   438 => x"06863883",
   439 => x"ffe1a054",
   440 => x"7281df06",
   441 => x"f0057081",
   442 => x"ff065153",
   443 => x"b8732789",
   444 => x"38ef1370",
   445 => x"81ff0651",
   446 => x"5374842b",
   447 => x"730755a0",
   448 => x"808d9604",
   449 => x"72a32ea1",
   450 => x"38737081",
   451 => x"0555a080",
   452 => x"80ae2d53",
   453 => x"72a02ef1",
   454 => x"38ff1475",
   455 => x"53705254",
   456 => x"a0809ba8",
   457 => x"2d74fc80",
   458 => x"0c737081",
   459 => x"0555a080",
   460 => x"80ae2d53",
   461 => x"728a2e09",
   462 => x"8106ee38",
   463 => x"a0808d94",
   464 => x"04a0809f",
   465 => x"fc51a080",
   466 => x"83d92d80",
   467 => x"0b83ffe0",
   468 => x"800c0294",
   469 => x"050d0402",
   470 => x"e8050d77",
   471 => x"797b5855",
   472 => x"55805372",
   473 => x"7625ab38",
   474 => x"74708105",
   475 => x"56a08080",
   476 => x"ae2d7470",
   477 => x"810556a0",
   478 => x"8080ae2d",
   479 => x"52527171",
   480 => x"2e883881",
   481 => x"51a0808f",
   482 => x"94048113",
   483 => x"53a0808e",
   484 => x"e3048051",
   485 => x"7083ffe0",
   486 => x"800c0298",
   487 => x"050d0402",
   488 => x"d8050dff",
   489 => x"0b83fff5",
   490 => x"cc0c800b",
   491 => x"83fff5e0",
   492 => x"0ca080a0",
   493 => x"8851a080",
   494 => x"83d92d83",
   495 => x"fff1b852",
   496 => x"8051a080",
   497 => x"8aa02d83",
   498 => x"ffe08008",
   499 => x"5483ffe0",
   500 => x"80089238",
   501 => x"a080a098",
   502 => x"51a08083",
   503 => x"d92d7355",
   504 => x"a0809783",
   505 => x"04a080a0",
   506 => x"ac51a080",
   507 => x"83d92d80",
   508 => x"56810b83",
   509 => x"fff1ac0c",
   510 => x"8853a080",
   511 => x"a0c45283",
   512 => x"fff1ee51",
   513 => x"a0808ed7",
   514 => x"2d83ffe0",
   515 => x"8008762e",
   516 => x"0981068b",
   517 => x"3883ffe0",
   518 => x"800883ff",
   519 => x"f1ac0c88",
   520 => x"53a080a0",
   521 => x"d05283ff",
   522 => x"f28a51a0",
   523 => x"808ed72d",
   524 => x"83ffe080",
   525 => x"088b3883",
   526 => x"ffe08008",
   527 => x"83fff1ac",
   528 => x"0c83fff1",
   529 => x"ac0852a0",
   530 => x"80a0dc51",
   531 => x"a0808181",
   532 => x"2d83fff1",
   533 => x"ac08802e",
   534 => x"81bb3883",
   535 => x"fff4fe0b",
   536 => x"a08080ae",
   537 => x"2d83fff4",
   538 => x"ff0ba080",
   539 => x"80ae2d71",
   540 => x"982b7190",
   541 => x"2b0783ff",
   542 => x"f5800ba0",
   543 => x"8080ae2d",
   544 => x"70882b72",
   545 => x"0783fff5",
   546 => x"810ba080",
   547 => x"80ae2d71",
   548 => x"0783fff5",
   549 => x"b60ba080",
   550 => x"80ae2d83",
   551 => x"fff5b70b",
   552 => x"a08080ae",
   553 => x"2d71882b",
   554 => x"07535f54",
   555 => x"525a5657",
   556 => x"557381ab",
   557 => x"aa2e0981",
   558 => x"06933875",
   559 => x"51a0808b",
   560 => x"cf2d83ff",
   561 => x"e0800856",
   562 => x"a08091e3",
   563 => x"047382d4",
   564 => x"d52e9038",
   565 => x"a080a0f0",
   566 => x"51a08083",
   567 => x"d92da080",
   568 => x"93db0475",
   569 => x"52a080a1",
   570 => x"9051a080",
   571 => x"81812d83",
   572 => x"fff1b852",
   573 => x"7551a080",
   574 => x"8aa02d83",
   575 => x"ffe08008",
   576 => x"5583ffe0",
   577 => x"8008802e",
   578 => x"84f938a0",
   579 => x"80a1a851",
   580 => x"a08083d9",
   581 => x"2da080a1",
   582 => x"d051a080",
   583 => x"81812d88",
   584 => x"53a080a0",
   585 => x"d05283ff",
   586 => x"f28a51a0",
   587 => x"808ed72d",
   588 => x"83ffe080",
   589 => x"088d3881",
   590 => x"0b83fff5",
   591 => x"e00ca080",
   592 => x"92ec0488",
   593 => x"53a080a0",
   594 => x"c45283ff",
   595 => x"f1ee51a0",
   596 => x"808ed72d",
   597 => x"83ffe080",
   598 => x"08802e90",
   599 => x"38a080a1",
   600 => x"e851a080",
   601 => x"81812da0",
   602 => x"8093db04",
   603 => x"83fff5b6",
   604 => x"0ba08080",
   605 => x"ae2d5473",
   606 => x"80d52e09",
   607 => x"810680db",
   608 => x"3883fff5",
   609 => x"b70ba080",
   610 => x"80ae2d54",
   611 => x"7381aa2e",
   612 => x"09810680",
   613 => x"c638800b",
   614 => x"83fff1b8",
   615 => x"0ba08080",
   616 => x"ae2d5654",
   617 => x"7481e92e",
   618 => x"83388154",
   619 => x"7481eb2e",
   620 => x"8c388055",
   621 => x"73752e09",
   622 => x"810683c7",
   623 => x"3883fff1",
   624 => x"c30ba080",
   625 => x"80ae2d55",
   626 => x"74913883",
   627 => x"fff1c40b",
   628 => x"a08080ae",
   629 => x"2d547382",
   630 => x"2e883880",
   631 => x"55a08097",
   632 => x"830483ff",
   633 => x"f1c50ba0",
   634 => x"8080ae2d",
   635 => x"7083fff5",
   636 => x"e80cff05",
   637 => x"83fff5dc",
   638 => x"0c83fff1",
   639 => x"c60ba080",
   640 => x"80ae2d83",
   641 => x"fff1c70b",
   642 => x"a08080ae",
   643 => x"2d587605",
   644 => x"77828029",
   645 => x"057083ff",
   646 => x"f5d00c83",
   647 => x"fff1c80b",
   648 => x"a08080ae",
   649 => x"2d7083ff",
   650 => x"f5c80c83",
   651 => x"fff5e008",
   652 => x"59575876",
   653 => x"802e81df",
   654 => x"388853a0",
   655 => x"80a0d052",
   656 => x"83fff28a",
   657 => x"51a0808e",
   658 => x"d72d83ff",
   659 => x"e0800882",
   660 => x"b23883ff",
   661 => x"f5e80870",
   662 => x"842b83ff",
   663 => x"f5b80c70",
   664 => x"83fff5e4",
   665 => x"0c83fff1",
   666 => x"dd0ba080",
   667 => x"80ae2d83",
   668 => x"fff1dc0b",
   669 => x"a08080ae",
   670 => x"2d718280",
   671 => x"290583ff",
   672 => x"f1de0ba0",
   673 => x"8080ae2d",
   674 => x"70848080",
   675 => x"291283ff",
   676 => x"f1df0ba0",
   677 => x"8080ae2d",
   678 => x"7081800a",
   679 => x"29127083",
   680 => x"fff1b00c",
   681 => x"83fff5c8",
   682 => x"08712983",
   683 => x"fff5d008",
   684 => x"057083ff",
   685 => x"f5f00c83",
   686 => x"fff1e50b",
   687 => x"a08080ae",
   688 => x"2d83fff1",
   689 => x"e40ba080",
   690 => x"80ae2d71",
   691 => x"82802905",
   692 => x"83fff1e6",
   693 => x"0ba08080",
   694 => x"ae2d7084",
   695 => x"80802912",
   696 => x"83fff1e7",
   697 => x"0ba08080",
   698 => x"ae2d7098",
   699 => x"2b81f00a",
   700 => x"06720570",
   701 => x"83fff1b4",
   702 => x"0cfe117e",
   703 => x"29770583",
   704 => x"fff5d80c",
   705 => x"52595243",
   706 => x"545e5152",
   707 => x"59525d57",
   708 => x"5957a080",
   709 => x"97810483",
   710 => x"fff1ca0b",
   711 => x"a08080ae",
   712 => x"2d83fff1",
   713 => x"c90ba080",
   714 => x"80ae2d71",
   715 => x"82802905",
   716 => x"7083fff5",
   717 => x"b80c70a0",
   718 => x"2983ff05",
   719 => x"70892a70",
   720 => x"83fff5e4",
   721 => x"0c83fff1",
   722 => x"cf0ba080",
   723 => x"80ae2d83",
   724 => x"fff1ce0b",
   725 => x"a08080ae",
   726 => x"2d718280",
   727 => x"29057083",
   728 => x"fff1b00c",
   729 => x"7b71291e",
   730 => x"7083fff5",
   731 => x"d80c7d83",
   732 => x"fff1b40c",
   733 => x"730583ff",
   734 => x"f5f00c55",
   735 => x"5e515155",
   736 => x"55815574",
   737 => x"83ffe080",
   738 => x"0c02a805",
   739 => x"0d0402ec",
   740 => x"050d7670",
   741 => x"872c7180",
   742 => x"ff065755",
   743 => x"5383fff5",
   744 => x"e0088a38",
   745 => x"72882c73",
   746 => x"81ff0656",
   747 => x"547383ff",
   748 => x"f5cc082e",
   749 => x"a83883ff",
   750 => x"f1b85283",
   751 => x"fff5d008",
   752 => x"1451a080",
   753 => x"8aa02d83",
   754 => x"ffe08008",
   755 => x"5383ffe0",
   756 => x"8008802e",
   757 => x"80cb3873",
   758 => x"83fff5cc",
   759 => x"0c83fff5",
   760 => x"e008802e",
   761 => x"a0387484",
   762 => x"2983fff1",
   763 => x"b8057008",
   764 => x"5253a080",
   765 => x"8bcf2d83",
   766 => x"ffe08008",
   767 => x"f00a0655",
   768 => x"a080989f",
   769 => x"04741083",
   770 => x"fff1b805",
   771 => x"70a08080",
   772 => x"992d5253",
   773 => x"a0808c81",
   774 => x"2d83ffe0",
   775 => x"80085574",
   776 => x"537283ff",
   777 => x"e0800c02",
   778 => x"94050d04",
   779 => x"02cc050d",
   780 => x"7e605e5b",
   781 => x"8056ff0b",
   782 => x"83fff5cc",
   783 => x"0c83fff1",
   784 => x"b40883ff",
   785 => x"f5d80856",
   786 => x"5783fff5",
   787 => x"e008762e",
   788 => x"8e3883ff",
   789 => x"f5e80884",
   790 => x"2b59a080",
   791 => x"98e70483",
   792 => x"fff5e408",
   793 => x"842b5980",
   794 => x"5a797927",
   795 => x"81e13879",
   796 => x"8f06a017",
   797 => x"575473a1",
   798 => x"387452a0",
   799 => x"80a28851",
   800 => x"a0808181",
   801 => x"2d83fff1",
   802 => x"b8527451",
   803 => x"811555a0",
   804 => x"808aa02d",
   805 => x"83fff1b8",
   806 => x"568076a0",
   807 => x"8080ae2d",
   808 => x"55587378",
   809 => x"2e833881",
   810 => x"587381e5",
   811 => x"2e819838",
   812 => x"81707906",
   813 => x"555c7380",
   814 => x"2e818c38",
   815 => x"8b16a080",
   816 => x"80ae2d98",
   817 => x"06587780",
   818 => x"fe388b53",
   819 => x"7c527551",
   820 => x"a0808ed7",
   821 => x"2d83ffe0",
   822 => x"800880eb",
   823 => x"389c1608",
   824 => x"51a0808b",
   825 => x"cf2d83ff",
   826 => x"e0800884",
   827 => x"1c0c9a16",
   828 => x"a0808099",
   829 => x"2d51a080",
   830 => x"8c812d83",
   831 => x"ffe08008",
   832 => x"83ffe080",
   833 => x"08555583",
   834 => x"fff5e008",
   835 => x"802e9e38",
   836 => x"9416a080",
   837 => x"80992d51",
   838 => x"a0808c81",
   839 => x"2d83ffe0",
   840 => x"8008902b",
   841 => x"83fff00a",
   842 => x"06701651",
   843 => x"5473881c",
   844 => x"0c777b0c",
   845 => x"7c52a080",
   846 => x"a2a851a0",
   847 => x"8081812d",
   848 => x"7b54a080",
   849 => x"9b9d0481",
   850 => x"1a5aa080",
   851 => x"98e90483",
   852 => x"fff5e008",
   853 => x"802e80c3",
   854 => x"387651a0",
   855 => x"80978e2d",
   856 => x"83ffe080",
   857 => x"0883ffe0",
   858 => x"800853a0",
   859 => x"80a2bc52",
   860 => x"57a08081",
   861 => x"812d7680",
   862 => x"fffffff8",
   863 => x"06547380",
   864 => x"fffffff8",
   865 => x"2e9538fe",
   866 => x"1783fff5",
   867 => x"e8082983",
   868 => x"fff5f008",
   869 => x"0555a080",
   870 => x"98e70480",
   871 => x"547383ff",
   872 => x"e0800c02",
   873 => x"b4050d04",
   874 => x"02e4050d",
   875 => x"787a7154",
   876 => x"83fff5bc",
   877 => x"535555a0",
   878 => x"8098ac2d",
   879 => x"83ffe080",
   880 => x"0881ff06",
   881 => x"5372802e",
   882 => x"818338a0",
   883 => x"80a2d451",
   884 => x"a08083d9",
   885 => x"2d83fff5",
   886 => x"c00883ff",
   887 => x"05892a57",
   888 => x"80705656",
   889 => x"75772581",
   890 => x"803883ff",
   891 => x"f5c408fe",
   892 => x"0583fff5",
   893 => x"e8082983",
   894 => x"fff5f008",
   895 => x"117683ff",
   896 => x"f5dc0806",
   897 => x"05755452",
   898 => x"53a0808a",
   899 => x"a02d83ff",
   900 => x"e0800880",
   901 => x"2e80c738",
   902 => x"81157083",
   903 => x"fff5dc08",
   904 => x"06545572",
   905 => x"963883ff",
   906 => x"f5c40851",
   907 => x"a080978e",
   908 => x"2d83ffe0",
   909 => x"800883ff",
   910 => x"f5c40c84",
   911 => x"80148117",
   912 => x"57547676",
   913 => x"24ffa338",
   914 => x"a0809ce9",
   915 => x"047452a0",
   916 => x"80a2f051",
   917 => x"a0808181",
   918 => x"2da0809c",
   919 => x"eb0483ff",
   920 => x"e0800853",
   921 => x"a0809ceb",
   922 => x"04815372",
   923 => x"83ffe080",
   924 => x"0c029c05",
   925 => x"0d0483ff",
   926 => x"e08c0802",
   927 => x"83ffe08c",
   928 => x"0cff3d0d",
   929 => x"800b83ff",
   930 => x"e08c08fc",
   931 => x"050c83ff",
   932 => x"e08c0888",
   933 => x"05088106",
   934 => x"ff117009",
   935 => x"7083ffe0",
   936 => x"8c088c05",
   937 => x"080683ff",
   938 => x"e08c08fc",
   939 => x"05081183",
   940 => x"ffe08c08",
   941 => x"fc050c83",
   942 => x"ffe08c08",
   943 => x"88050881",
   944 => x"2a83ffe0",
   945 => x"8c088805",
   946 => x"0c83ffe0",
   947 => x"8c088c05",
   948 => x"081083ff",
   949 => x"e08c088c",
   950 => x"050c5151",
   951 => x"515183ff",
   952 => x"e08c0888",
   953 => x"0508802e",
   954 => x"8438ffa2",
   955 => x"3983ffe0",
   956 => x"8c08fc05",
   957 => x"087083ff",
   958 => x"e0800c51",
   959 => x"833d0d83",
   960 => x"ffe08c0c",
   961 => x"04000000",
   962 => x"00ffffff",
   963 => x"ff00ffff",
   964 => x"ffff00ff",
   965 => x"ffffff00",
   966 => x"436d645f",
   967 => x"696e6974",
   968 => x"0a000000",
   969 => x"636d645f",
   970 => x"434d4438",
   971 => x"20726573",
   972 => x"706f6e73",
   973 => x"653a2025",
   974 => x"640a0000",
   975 => x"53444843",
   976 => x"20496e69",
   977 => x"7469616c",
   978 => x"697a6174",
   979 => x"696f6e20",
   980 => x"6572726f",
   981 => x"72210a00",
   982 => x"434d4438",
   983 => x"5f342072",
   984 => x"6573706f",
   985 => x"6e73653a",
   986 => x"2025640a",
   987 => x"00000000",
   988 => x"434d4435",
   989 => x"38202564",
   990 => x"0a202000",
   991 => x"434d4435",
   992 => x"385f3220",
   993 => x"25640a20",
   994 => x"20000000",
   995 => x"52656164",
   996 => x"20636f6d",
   997 => x"6d616e64",
   998 => x"20666169",
   999 => x"6c656420",
  1000 => x"61742025",
  1001 => x"64202825",
  1002 => x"64290a00",
  1003 => x"496e6974",
  1004 => x"69616c69",
  1005 => x"7a696e67",
  1006 => x"20534420",
  1007 => x"63617264",
  1008 => x"0a000000",
  1009 => x"48756e74",
  1010 => x"696e6720",
  1011 => x"666f7220",
  1012 => x"70617274",
  1013 => x"6974696f",
  1014 => x"6e0a0000",
  1015 => x"4d414e49",
  1016 => x"46455354",
  1017 => x"4d535400",
  1018 => x"50617273",
  1019 => x"696e6720",
  1020 => x"6d616e69",
  1021 => x"66657374",
  1022 => x"0a000000",
  1023 => x"52657475",
  1024 => x"726e696e",
  1025 => x"670a0000",
  1026 => x"52656164",
  1027 => x"696e6720",
  1028 => x"4d42520a",
  1029 => x"00000000",
  1030 => x"52656164",
  1031 => x"206f6620",
  1032 => x"4d425220",
  1033 => x"6661696c",
  1034 => x"65640a00",
  1035 => x"4d425220",
  1036 => x"73756363",
  1037 => x"65737366",
  1038 => x"756c6c79",
  1039 => x"20726561",
  1040 => x"640a0000",
  1041 => x"46415431",
  1042 => x"36202020",
  1043 => x"00000000",
  1044 => x"46415433",
  1045 => x"32202020",
  1046 => x"00000000",
  1047 => x"50617274",
  1048 => x"6974696f",
  1049 => x"6e636f75",
  1050 => x"6e742025",
  1051 => x"640a0000",
  1052 => x"4e6f2070",
  1053 => x"61727469",
  1054 => x"74696f6e",
  1055 => x"20736967",
  1056 => x"6e617475",
  1057 => x"72652066",
  1058 => x"6f756e64",
  1059 => x"0a000000",
  1060 => x"52656164",
  1061 => x"696e6720",
  1062 => x"626f6f74",
  1063 => x"20736563",
  1064 => x"746f7220",
  1065 => x"25640a00",
  1066 => x"52656164",
  1067 => x"20626f6f",
  1068 => x"74207365",
  1069 => x"63746f72",
  1070 => x"2066726f",
  1071 => x"6d206669",
  1072 => x"72737420",
  1073 => x"70617274",
  1074 => x"6974696f",
  1075 => x"6e0a0000",
  1076 => x"48756e74",
  1077 => x"696e6720",
  1078 => x"666f7220",
  1079 => x"66696c65",
  1080 => x"73797374",
  1081 => x"656d0a00",
  1082 => x"556e7375",
  1083 => x"70706f72",
  1084 => x"74656420",
  1085 => x"70617274",
  1086 => x"6974696f",
  1087 => x"6e207479",
  1088 => x"7065210d",
  1089 => x"00000000",
  1090 => x"52656164",
  1091 => x"696e6720",
  1092 => x"64697265",
  1093 => x"63746f72",
  1094 => x"79207365",
  1095 => x"63746f72",
  1096 => x"2025640a",
  1097 => x"00000000",
  1098 => x"66696c65",
  1099 => x"20222573",
  1100 => x"2220666f",
  1101 => x"756e640d",
  1102 => x"00000000",
  1103 => x"47657446",
  1104 => x"41544c69",
  1105 => x"6e6b2072",
  1106 => x"65747572",
  1107 => x"6e656420",
  1108 => x"25640a00",
  1109 => x"4f70656e",
  1110 => x"65642066",
  1111 => x"696c652c",
  1112 => x"206c6f61",
  1113 => x"64696e67",
  1114 => x"2e2e2e0a",
  1115 => x"00000000",
  1116 => x"43616e27",
  1117 => x"74206f70",
  1118 => x"656e2025",
  1119 => x"730a0000",
	others => x"00000000"
);

begin

process (clk)
begin
	if (clk'event and clk = '1') then
		if (from_zpu.memAWriteEnable = '1') and (from_zpu.memBWriteEnable = '1') and (from_zpu.memAAddr=from_zpu.memBAddr) and (from_zpu.memAWrite/=from_zpu.memBWrite) then
			report "write collision" severity failure;
		end if;
	
		if (from_zpu.memAWriteEnable = '1') then
			ram(to_integer(unsigned(from_zpu.memAAddr(maxAddrBitBRAM downto 2)))) := from_zpu.memAWrite;
			to_zpu.memARead <= from_zpu.memAWrite;
		else
			to_zpu.memARead <= ram(to_integer(unsigned(from_zpu.memAAddr(maxAddrBitBRAM downto 2))));
		end if;
	end if;
end process;

process (clk)
begin
	if (clk'event and clk = '1') then
		if (from_zpu.memBWriteEnable = '1') then
			ram(to_integer(unsigned(from_zpu.memBAddr(maxAddrBitBRAM downto 2)))) := from_zpu.memBWrite;
			to_zpu.memBRead <= from_zpu.memBWrite;
		else
			to_zpu.memBRead <= ram(to_integer(unsigned(from_zpu.memBAddr(maxAddrBitBRAM downto 2))));
		end if;
	end if;
end process;


end arch;

