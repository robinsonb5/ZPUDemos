-- ZPU
--
-- Copyright 2004-2008 oharboe - �yvind Harboe - oyvind.harboe@zylin.com
-- Modified by Alastair M. Robinson for the ZPUFlex project.
--
-- The FreeBSD license
-- 
-- Redistribution and use in source and binary forms, with or without
-- modification, are permitted provided that the following conditions
-- are met:
-- 
-- 1. Redistributions of source code must retain the above copyright
--    notice, this list of conditions and the following disclaimer.
-- 2. Redistributions in binary form must reproduce the above
--    copyright notice, this list of conditions and the following
--    disclaimer in the documentation and/or other materials
--    provided with the distribution.
-- 
-- THIS SOFTWARE IS PROVIDED BY THE ZPU PROJECT ``AS IS'' AND ANY
-- EXPRESS OR IMPLIED WARRANTIES, INCLUDING, BUT NOT LIMITED TO,
-- THE IMPLIED WARRANTIES OF MERCHANTABILITY AND FITNESS FOR A
-- PARTICULAR PURPOSE ARE DISCLAIMED. IN NO EVENT SHALL THE
-- ZPU PROJECT OR CONTRIBUTORS BE LIABLE FOR ANY DIRECT,
-- INDIRECT, INCIDENTAL, SPECIAL, EXEMPLARY, OR CONSEQUENTIAL DAMAGES
-- (INCLUDING, BUT NOT LIMITED TO, PROCUREMENT OF SUBSTITUTE GOODS
-- OR SERVICES; LOSS OF USE, DATA, OR PROFITS; OR BUSINESS INTERRUPTION)
-- HOWEVER CAUSED AND ON ANY THEORY OF LIABILITY, WHETHER IN CONTRACT,
-- STRICT LIABILITY, OR TORT (INCLUDING NEGLIGENCE OR OTHERWISE)
-- ARISING IN ANY WAY OUT OF THE USE OF THIS SOFTWARE, EVEN IF
-- ADVISED OF THE POSSIBILITY OF SUCH DAMAGE.
-- 
-- The views and conclusions contained in the software and documentation
-- are those of the authors and should not be interpreted as representing
-- official policies, either expressed or implied, of the ZPU Project.

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;


library work;
use work.zpu_config.all;
use work.zpupkg.all;

entity SDBootstrap_ROM is
generic
	(
		maxAddrBitBRAM : integer := maxAddrBitBRAMLimit -- Specify your actual ROM size to save LEs and unnecessary block RAM usage.
	);
port (
	clk : in std_logic;
	areset : in std_logic := '0';
	from_zpu : in ZPU_ToROM;
	to_zpu : out ZPU_FromROM
);
end SDBootstrap_ROM;

architecture arch of SDBootstrap_ROM is

type ram_type is array(natural range 0 to ((2**(maxAddrBitBRAM+1))/4)-1) of std_logic_vector(wordSize-1 downto 0);

shared variable ram : ram_type :=
(
     0 => x"84808080",
     1 => x"ed040000",
     2 => x"00000000",
     3 => x"84808080",
     4 => x"880d8004",
     5 => x"84808080",
     6 => x"940471fd",
     7 => x"06087283",
     8 => x"06098105",
     9 => x"8205832b",
    10 => x"2a83ffff",
    11 => x"06520471",
    12 => x"fc060872",
    13 => x"83060981",
    14 => x"05830510",
    15 => x"10102a81",
    16 => x"ff065204",
    17 => x"71fc0608",
    18 => x"8480809f",
    19 => x"e8738306",
    20 => x"10100508",
    21 => x"067381ff",
    22 => x"06738306",
    23 => x"09810583",
    24 => x"05101010",
    25 => x"2b0772fc",
    26 => x"060c5151",
    27 => x"04028405",
    28 => x"84808080",
    29 => x"880c8480",
    30 => x"8080940b",
    31 => x"8480808d",
    32 => x"9d040000",
    33 => x"02c4050d",
    34 => x"0280c005",
    35 => x"83ffe0e0",
    36 => x"5b568076",
    37 => x"70840558",
    38 => x"08715e5e",
    39 => x"577c7084",
    40 => x"055e0858",
    41 => x"805b7798",
    42 => x"2a78882b",
    43 => x"59547389",
    44 => x"38765e84",
    45 => x"808083e3",
    46 => x"047b802e",
    47 => x"81fd3880",
    48 => x"5c7380e4",
    49 => x"2ea13873",
    50 => x"80e4268e",
    51 => x"387380e3",
    52 => x"2e819a38",
    53 => x"84808082",
    54 => x"fb047380",
    55 => x"f32e80f5",
    56 => x"38848080",
    57 => x"82fb0475",
    58 => x"84177108",
    59 => x"7e5c5557",
    60 => x"52728025",
    61 => x"8e38ad51",
    62 => x"84808083",
    63 => x"ee2d7209",
    64 => x"81055372",
    65 => x"802ebe38",
    66 => x"8755729c",
    67 => x"2a73842b",
    68 => x"54527180",
    69 => x"2e833881",
    70 => x"59897225",
    71 => x"8a38b712",
    72 => x"52848080",
    73 => x"82aa04b0",
    74 => x"12527880",
    75 => x"2e893871",
    76 => x"51848080",
    77 => x"83ee2dff",
    78 => x"15557480",
    79 => x"25cc3884",
    80 => x"808082cd",
    81 => x"04b05184",
    82 => x"808083ee",
    83 => x"2d805384",
    84 => x"80808394",
    85 => x"04758417",
    86 => x"71087054",
    87 => x"5c575284",
    88 => x"80808492",
    89 => x"2d7b5384",
    90 => x"80808394",
    91 => x"04758417",
    92 => x"71085657",
    93 => x"52848080",
    94 => x"83cb04a5",
    95 => x"51848080",
    96 => x"83ee2d73",
    97 => x"51848080",
    98 => x"83ee2d82",
    99 => x"17578480",
   100 => x"8083d604",
   101 => x"72ff1454",
   102 => x"52807225",
   103 => x"b9387970",
   104 => x"81055b84",
   105 => x"808080af",
   106 => x"2d705254",
   107 => x"84808083",
   108 => x"ee2d8117",
   109 => x"57848080",
   110 => x"83940473",
   111 => x"a52e0981",
   112 => x"06893881",
   113 => x"5c848080",
   114 => x"83d60473",
   115 => x"51848080",
   116 => x"83ee2d81",
   117 => x"1757811b",
   118 => x"5b837b25",
   119 => x"fdc83873",
   120 => x"fdbb387d",
   121 => x"83ffe080",
   122 => x"0c02bc05",
   123 => x"0d0402f8",
   124 => x"050d7352",
   125 => x"c0087088",
   126 => x"2a708106",
   127 => x"51515170",
   128 => x"802ef138",
   129 => x"71c00c71",
   130 => x"83ffe080",
   131 => x"0c028805",
   132 => x"0d0402e8",
   133 => x"050d8078",
   134 => x"57557570",
   135 => x"84055708",
   136 => x"53805472",
   137 => x"982a7388",
   138 => x"2b545271",
   139 => x"802ea238",
   140 => x"c0087088",
   141 => x"2a708106",
   142 => x"51515170",
   143 => x"802ef138",
   144 => x"71c00c81",
   145 => x"15811555",
   146 => x"55837425",
   147 => x"d63871ca",
   148 => x"387483ff",
   149 => x"e0800c02",
   150 => x"98050d04",
   151 => x"02f4050d",
   152 => x"74767181",
   153 => x"ff06d40c",
   154 => x"535383ff",
   155 => x"f1a00885",
   156 => x"3871892b",
   157 => x"5271982a",
   158 => x"d40c7190",
   159 => x"2a7081ff",
   160 => x"06d40c51",
   161 => x"71882a70",
   162 => x"81ff06d4",
   163 => x"0c517181",
   164 => x"ff06d40c",
   165 => x"72902a70",
   166 => x"81ff06d4",
   167 => x"0c51d408",
   168 => x"7081ff06",
   169 => x"515182b8",
   170 => x"bf527081",
   171 => x"ff2e0981",
   172 => x"06943881",
   173 => x"ff0bd40c",
   174 => x"d4087081",
   175 => x"ff06ff14",
   176 => x"54515171",
   177 => x"e5387083",
   178 => x"ffe0800c",
   179 => x"028c050d",
   180 => x"0402fc05",
   181 => x"0d81c751",
   182 => x"81ff0bd4",
   183 => x"0cff1151",
   184 => x"708025f4",
   185 => x"38028405",
   186 => x"0d0402f0",
   187 => x"050d8480",
   188 => x"8085d12d",
   189 => x"819c9f53",
   190 => x"805287fc",
   191 => x"80f75184",
   192 => x"808084dc",
   193 => x"2d83ffe0",
   194 => x"80085483",
   195 => x"ffe08008",
   196 => x"812e0981",
   197 => x"06ae3881",
   198 => x"ff0bd40c",
   199 => x"820a5284",
   200 => x"9c80e951",
   201 => x"84808084",
   202 => x"dc2d83ff",
   203 => x"e080088e",
   204 => x"3881ff0b",
   205 => x"d40c7353",
   206 => x"84808086",
   207 => x"cb048480",
   208 => x"8085d12d",
   209 => x"ff135372",
   210 => x"ffae3872",
   211 => x"83ffe080",
   212 => x"0c029005",
   213 => x"0d0402f4",
   214 => x"050d81ff",
   215 => x"0bd40c84",
   216 => x"80809ff8",
   217 => x"51848080",
   218 => x"84922d93",
   219 => x"53805287",
   220 => x"fc80c151",
   221 => x"84808084",
   222 => x"dc2d83ff",
   223 => x"e080088e",
   224 => x"3881ff0b",
   225 => x"d40c8153",
   226 => x"84808087",
   227 => x"9a048480",
   228 => x"8085d12d",
   229 => x"ff135372",
   230 => x"d4387283",
   231 => x"ffe0800c",
   232 => x"028c050d",
   233 => x"0402f005",
   234 => x"0d848080",
   235 => x"85d12d83",
   236 => x"aa52849c",
   237 => x"80c85184",
   238 => x"808084dc",
   239 => x"2d83ffe0",
   240 => x"800883ff",
   241 => x"e0800853",
   242 => x"848080a0",
   243 => x"84525484",
   244 => x"80808184",
   245 => x"2d73812e",
   246 => x"09810690",
   247 => x"38d80870",
   248 => x"83ffff06",
   249 => x"54547283",
   250 => x"aa2ea938",
   251 => x"84808086",
   252 => x"d62d8480",
   253 => x"80888c04",
   254 => x"81548480",
   255 => x"8089c304",
   256 => x"848080a0",
   257 => x"9c518480",
   258 => x"8081842d",
   259 => x"80548480",
   260 => x"8089c304",
   261 => x"73528480",
   262 => x"80a0b851",
   263 => x"84808081",
   264 => x"842d81ff",
   265 => x"0bd40cb1",
   266 => x"53848080",
   267 => x"85ea2d83",
   268 => x"ffe08008",
   269 => x"802e80fc",
   270 => x"38805287",
   271 => x"fc80fa51",
   272 => x"84808084",
   273 => x"dc2d83ff",
   274 => x"e0800880",
   275 => x"d53883ff",
   276 => x"e0800852",
   277 => x"848080a0",
   278 => x"d0518480",
   279 => x"8081842d",
   280 => x"81ff0bd4",
   281 => x"0cd40881",
   282 => x"ff067053",
   283 => x"848080a0",
   284 => x"dc525484",
   285 => x"80808184",
   286 => x"2d81ff0b",
   287 => x"d40c81ff",
   288 => x"0bd40c81",
   289 => x"ff0bd40c",
   290 => x"81ff0bd4",
   291 => x"0c73862a",
   292 => x"70810670",
   293 => x"56515372",
   294 => x"802ea838",
   295 => x"84808087",
   296 => x"f80483ff",
   297 => x"e0800852",
   298 => x"848080a0",
   299 => x"d0518480",
   300 => x"8081842d",
   301 => x"72822efe",
   302 => x"c738ff13",
   303 => x"5372fee9",
   304 => x"38725473",
   305 => x"83ffe080",
   306 => x"0c029005",
   307 => x"0d0402f4",
   308 => x"050d810b",
   309 => x"83fff1a0",
   310 => x"0cd00870",
   311 => x"8f2a7081",
   312 => x"06515153",
   313 => x"72f33872",
   314 => x"d00c8480",
   315 => x"8085d12d",
   316 => x"d008708f",
   317 => x"2a708106",
   318 => x"51515372",
   319 => x"f338810b",
   320 => x"d00c8753",
   321 => x"805284d4",
   322 => x"80c05184",
   323 => x"808084dc",
   324 => x"2d83ffe0",
   325 => x"8008812e",
   326 => x"97387282",
   327 => x"2e098106",
   328 => x"89388053",
   329 => x"8480808a",
   330 => x"ea04ff13",
   331 => x"5372d538",
   332 => x"84808087",
   333 => x"a52d83ff",
   334 => x"e0800883",
   335 => x"fff1a00c",
   336 => x"815287fc",
   337 => x"80d05184",
   338 => x"808084dc",
   339 => x"2d81ff0b",
   340 => x"d40cd008",
   341 => x"708f2a70",
   342 => x"81065151",
   343 => x"5372f338",
   344 => x"72d00c81",
   345 => x"ff0bd40c",
   346 => x"81537283",
   347 => x"ffe0800c",
   348 => x"028c050d",
   349 => x"04800b83",
   350 => x"ffe0800c",
   351 => x"0402e005",
   352 => x"0d797b57",
   353 => x"57805881",
   354 => x"ff0bd40c",
   355 => x"d008708f",
   356 => x"2a708106",
   357 => x"51515473",
   358 => x"f3388281",
   359 => x"0bd00c81",
   360 => x"ff0bd40c",
   361 => x"765287fc",
   362 => x"80d15184",
   363 => x"808084dc",
   364 => x"2d80dbc6",
   365 => x"df5583ff",
   366 => x"e0800880",
   367 => x"2e9b3883",
   368 => x"ffe08008",
   369 => x"53765284",
   370 => x"8080a0ec",
   371 => x"51848080",
   372 => x"81842d84",
   373 => x"80808ca6",
   374 => x"0481ff0b",
   375 => x"d40cd408",
   376 => x"7081ff06",
   377 => x"51547381",
   378 => x"fe2e0981",
   379 => x"069c3880",
   380 => x"ff55d808",
   381 => x"76708405",
   382 => x"580cff15",
   383 => x"55748025",
   384 => x"f1388158",
   385 => x"8480808c",
   386 => x"9004ff15",
   387 => x"5574ca38",
   388 => x"81ff0bd4",
   389 => x"0cd00870",
   390 => x"8f2a7081",
   391 => x"06515154",
   392 => x"73f33873",
   393 => x"d00c7783",
   394 => x"ffe0800c",
   395 => x"02a0050d",
   396 => x"0402f405",
   397 => x"0d747088",
   398 => x"2a83fe80",
   399 => x"06707298",
   400 => x"2a077288",
   401 => x"2b87fc80",
   402 => x"80067398",
   403 => x"2b81f00a",
   404 => x"06717307",
   405 => x"0783ffe0",
   406 => x"800c5651",
   407 => x"5351028c",
   408 => x"050d0402",
   409 => x"f8050d02",
   410 => x"8e058480",
   411 => x"8080af2d",
   412 => x"74982b71",
   413 => x"902b0770",
   414 => x"902c83ff",
   415 => x"e0800c52",
   416 => x"52028805",
   417 => x"0d0402f8",
   418 => x"050d7370",
   419 => x"902b7190",
   420 => x"2a0783ff",
   421 => x"e0800c52",
   422 => x"0288050d",
   423 => x"0402ec05",
   424 => x"0d800bfc",
   425 => x"800c8480",
   426 => x"80a18c51",
   427 => x"84808084",
   428 => x"922d8480",
   429 => x"8089ce2d",
   430 => x"83ffe080",
   431 => x"08802e81",
   432 => x"f7388480",
   433 => x"80a1a451",
   434 => x"84808084",
   435 => x"922d8480",
   436 => x"80909c2d",
   437 => x"83ffe1a0",
   438 => x"52848080",
   439 => x"a1bc5184",
   440 => x"80809cff",
   441 => x"2d83ffe0",
   442 => x"8008802e",
   443 => x"81ca3883",
   444 => x"ffe1a00b",
   445 => x"848080a1",
   446 => x"c8525484",
   447 => x"80808492",
   448 => x"2d805573",
   449 => x"70810555",
   450 => x"84808080",
   451 => x"af2d5372",
   452 => x"a02e80e3",
   453 => x"3872a32e",
   454 => x"81843872",
   455 => x"80c72e09",
   456 => x"81068d38",
   457 => x"84808080",
   458 => x"8c2d8480",
   459 => x"808ed204",
   460 => x"728a2e09",
   461 => x"81068d38",
   462 => x"84808080",
   463 => x"942d8480",
   464 => x"808ed204",
   465 => x"7280cc2e",
   466 => x"09810686",
   467 => x"3883ffe1",
   468 => x"a0547281",
   469 => x"df06f005",
   470 => x"7081ff06",
   471 => x"5153b873",
   472 => x"278938ef",
   473 => x"137081ff",
   474 => x"06515374",
   475 => x"842b7307",
   476 => x"55848080",
   477 => x"8e830472",
   478 => x"a32ea338",
   479 => x"73708105",
   480 => x"55848080",
   481 => x"80af2d53",
   482 => x"72a02ef0",
   483 => x"38ff1475",
   484 => x"53705254",
   485 => x"8480809c",
   486 => x"ff2d74fc",
   487 => x"800c7370",
   488 => x"81055584",
   489 => x"808080af",
   490 => x"2d53728a",
   491 => x"2e098106",
   492 => x"ed388480",
   493 => x"808e8104",
   494 => x"848080a1",
   495 => x"dc518480",
   496 => x"8084922d",
   497 => x"800b83ff",
   498 => x"e0800c02",
   499 => x"94050d04",
   500 => x"02e8050d",
   501 => x"77797b58",
   502 => x"55558053",
   503 => x"727625af",
   504 => x"38747081",
   505 => x"05568480",
   506 => x"8080af2d",
   507 => x"74708105",
   508 => x"56848080",
   509 => x"80af2d52",
   510 => x"5271712e",
   511 => x"89388151",
   512 => x"84808090",
   513 => x"91048113",
   514 => x"53848080",
   515 => x"8fdc0480",
   516 => x"517083ff",
   517 => x"e0800c02",
   518 => x"98050d04",
   519 => x"02d8050d",
   520 => x"ff0b83ff",
   521 => x"f5cc0c80",
   522 => x"0b83fff5",
   523 => x"e00c8480",
   524 => x"80a1e851",
   525 => x"84808084",
   526 => x"922d83ff",
   527 => x"f1b85280",
   528 => x"51848080",
   529 => x"8afd2d83",
   530 => x"ffe08008",
   531 => x"5483ffe0",
   532 => x"80089538",
   533 => x"848080a1",
   534 => x"f8518480",
   535 => x"8084922d",
   536 => x"73558480",
   537 => x"8098c104",
   538 => x"848080a2",
   539 => x"8c518480",
   540 => x"8084922d",
   541 => x"8056810b",
   542 => x"83fff1ac",
   543 => x"0c885384",
   544 => x"8080a2a4",
   545 => x"5283fff1",
   546 => x"ee518480",
   547 => x"808fd02d",
   548 => x"83ffe080",
   549 => x"08762e09",
   550 => x"81068b38",
   551 => x"83ffe080",
   552 => x"0883fff1",
   553 => x"ac0c8853",
   554 => x"848080a2",
   555 => x"b05283ff",
   556 => x"f28a5184",
   557 => x"80808fd0",
   558 => x"2d83ffe0",
   559 => x"80088b38",
   560 => x"83ffe080",
   561 => x"0883fff1",
   562 => x"ac0c83ff",
   563 => x"f1ac0852",
   564 => x"848080a2",
   565 => x"bc518480",
   566 => x"8081842d",
   567 => x"83fff1ac",
   568 => x"08802e81",
   569 => x"cb3883ff",
   570 => x"f4fe0b84",
   571 => x"808080af",
   572 => x"2d83fff4",
   573 => x"ff0b8480",
   574 => x"8080af2d",
   575 => x"71982b71",
   576 => x"902b0783",
   577 => x"fff5800b",
   578 => x"84808080",
   579 => x"af2d7088",
   580 => x"2b720783",
   581 => x"fff5810b",
   582 => x"84808080",
   583 => x"af2d7107",
   584 => x"83fff5b6",
   585 => x"0b848080",
   586 => x"80af2d83",
   587 => x"fff5b70b",
   588 => x"84808080",
   589 => x"af2d7188",
   590 => x"2b07535f",
   591 => x"54525a56",
   592 => x"57557381",
   593 => x"abaa2e09",
   594 => x"81069538",
   595 => x"75518480",
   596 => x"808cb12d",
   597 => x"83ffe080",
   598 => x"08568480",
   599 => x"8092f904",
   600 => x"7382d4d5",
   601 => x"2e933884",
   602 => x"8080a2d0",
   603 => x"51848080",
   604 => x"84922d84",
   605 => x"80809585",
   606 => x"04755284",
   607 => x"8080a2f0",
   608 => x"51848080",
   609 => x"81842d83",
   610 => x"fff1b852",
   611 => x"75518480",
   612 => x"808afd2d",
   613 => x"83ffe080",
   614 => x"085583ff",
   615 => x"e0800880",
   616 => x"2e859e38",
   617 => x"848080a3",
   618 => x"88518480",
   619 => x"8084922d",
   620 => x"848080a3",
   621 => x"b0518480",
   622 => x"8081842d",
   623 => x"88538480",
   624 => x"80a2b052",
   625 => x"83fff28a",
   626 => x"51848080",
   627 => x"8fd02d83",
   628 => x"ffe08008",
   629 => x"8e38810b",
   630 => x"83fff5e0",
   631 => x"0c848080",
   632 => x"94910488",
   633 => x"53848080",
   634 => x"a2a45283",
   635 => x"fff1ee51",
   636 => x"8480808f",
   637 => x"d02d83ff",
   638 => x"e0800880",
   639 => x"2e933884",
   640 => x"8080a3c8",
   641 => x"51848080",
   642 => x"81842d84",
   643 => x"80809585",
   644 => x"0483fff5",
   645 => x"b60b8480",
   646 => x"8080af2d",
   647 => x"547380d5",
   648 => x"2e098106",
   649 => x"80df3883",
   650 => x"fff5b70b",
   651 => x"84808080",
   652 => x"af2d5473",
   653 => x"81aa2e09",
   654 => x"810680c9",
   655 => x"38800b83",
   656 => x"fff1b80b",
   657 => x"84808080",
   658 => x"af2d5654",
   659 => x"7481e92e",
   660 => x"83388154",
   661 => x"7481eb2e",
   662 => x"8c388055",
   663 => x"73752e09",
   664 => x"810683dd",
   665 => x"3883fff1",
   666 => x"c30b8480",
   667 => x"8080af2d",
   668 => x"55749238",
   669 => x"83fff1c4",
   670 => x"0b848080",
   671 => x"80af2d54",
   672 => x"73822e89",
   673 => x"38805584",
   674 => x"808098c1",
   675 => x"0483fff1",
   676 => x"c50b8480",
   677 => x"8080af2d",
   678 => x"7083fff5",
   679 => x"e80cff05",
   680 => x"83fff5dc",
   681 => x"0c83fff1",
   682 => x"c60b8480",
   683 => x"8080af2d",
   684 => x"83fff1c7",
   685 => x"0b848080",
   686 => x"80af2d58",
   687 => x"76057782",
   688 => x"80290570",
   689 => x"83fff5d0",
   690 => x"0c83fff1",
   691 => x"c80b8480",
   692 => x"8080af2d",
   693 => x"7083fff5",
   694 => x"c80c83ff",
   695 => x"f5e00859",
   696 => x"57587680",
   697 => x"2e81ea38",
   698 => x"88538480",
   699 => x"80a2b052",
   700 => x"83fff28a",
   701 => x"51848080",
   702 => x"8fd02d83",
   703 => x"ffe08008",
   704 => x"82bf3883",
   705 => x"fff5e808",
   706 => x"70842b83",
   707 => x"fff5b80c",
   708 => x"7083fff5",
   709 => x"e40c83ff",
   710 => x"f1dd0b84",
   711 => x"808080af",
   712 => x"2d83fff1",
   713 => x"dc0b8480",
   714 => x"8080af2d",
   715 => x"71828029",
   716 => x"0583fff1",
   717 => x"de0b8480",
   718 => x"8080af2d",
   719 => x"70848080",
   720 => x"291283ff",
   721 => x"f1df0b84",
   722 => x"808080af",
   723 => x"2d708180",
   724 => x"0a291270",
   725 => x"83fff1b0",
   726 => x"0c83fff5",
   727 => x"c8087129",
   728 => x"83fff5d0",
   729 => x"08057083",
   730 => x"fff5f00c",
   731 => x"83fff1e5",
   732 => x"0b848080",
   733 => x"80af2d83",
   734 => x"fff1e40b",
   735 => x"84808080",
   736 => x"af2d7182",
   737 => x"80290583",
   738 => x"fff1e60b",
   739 => x"84808080",
   740 => x"af2d7084",
   741 => x"80802912",
   742 => x"83fff1e7",
   743 => x"0b848080",
   744 => x"80af2d70",
   745 => x"982b81f0",
   746 => x"0a067205",
   747 => x"7083fff1",
   748 => x"b40cfe11",
   749 => x"7e297705",
   750 => x"83fff5d8",
   751 => x"0c525952",
   752 => x"43545e51",
   753 => x"5259525d",
   754 => x"57595784",
   755 => x"808098bf",
   756 => x"0483fff1",
   757 => x"ca0b8480",
   758 => x"8080af2d",
   759 => x"83fff1c9",
   760 => x"0b848080",
   761 => x"80af2d71",
   762 => x"82802905",
   763 => x"7083fff5",
   764 => x"b80c70a0",
   765 => x"2983ff05",
   766 => x"70892a70",
   767 => x"83fff5e4",
   768 => x"0c83fff1",
   769 => x"cf0b8480",
   770 => x"8080af2d",
   771 => x"83fff1ce",
   772 => x"0b848080",
   773 => x"80af2d71",
   774 => x"82802905",
   775 => x"7083fff1",
   776 => x"b00c7b71",
   777 => x"291e7083",
   778 => x"fff5d80c",
   779 => x"7d83fff1",
   780 => x"b40c7305",
   781 => x"83fff5f0",
   782 => x"0c555e51",
   783 => x"51555581",
   784 => x"557483ff",
   785 => x"e0800c02",
   786 => x"a8050d04",
   787 => x"02ec050d",
   788 => x"7670872c",
   789 => x"7180ff06",
   790 => x"57555383",
   791 => x"fff5e008",
   792 => x"8a387288",
   793 => x"2c7381ff",
   794 => x"06565473",
   795 => x"83fff5cc",
   796 => x"082ea938",
   797 => x"83fff1b8",
   798 => x"5283fff5",
   799 => x"d0081451",
   800 => x"8480808a",
   801 => x"fd2d83ff",
   802 => x"e0800853",
   803 => x"83ffe080",
   804 => x"08802e80",
   805 => x"cf387383",
   806 => x"fff5cc0c",
   807 => x"83fff5e0",
   808 => x"08802ea2",
   809 => x"38748429",
   810 => x"83fff1b8",
   811 => x"05700852",
   812 => x"53848080",
   813 => x"8cb12d83",
   814 => x"ffe08008",
   815 => x"f00a0655",
   816 => x"84808099",
   817 => x"e2047410",
   818 => x"83fff1b8",
   819 => x"05708480",
   820 => x"80809a2d",
   821 => x"52538480",
   822 => x"808ce32d",
   823 => x"83ffe080",
   824 => x"08557453",
   825 => x"7283ffe0",
   826 => x"800c0294",
   827 => x"050d0402",
   828 => x"cc050d7e",
   829 => x"605e5b80",
   830 => x"56ff0b83",
   831 => x"fff5cc0c",
   832 => x"83fff1b4",
   833 => x"0883fff5",
   834 => x"d8085657",
   835 => x"83fff5e0",
   836 => x"08762e8f",
   837 => x"3883fff5",
   838 => x"e808842b",
   839 => x"59848080",
   840 => x"9aab0483",
   841 => x"fff5e408",
   842 => x"842b5980",
   843 => x"5a797927",
   844 => x"81f03879",
   845 => x"8f06a017",
   846 => x"575473a4",
   847 => x"38745284",
   848 => x"8080a3e8",
   849 => x"51848080",
   850 => x"81842d83",
   851 => x"fff1b852",
   852 => x"74518115",
   853 => x"55848080",
   854 => x"8afd2d83",
   855 => x"fff1b856",
   856 => x"80768480",
   857 => x"8080af2d",
   858 => x"55587378",
   859 => x"2e833881",
   860 => x"587381e5",
   861 => x"2e81a238",
   862 => x"81707906",
   863 => x"555c7380",
   864 => x"2e819638",
   865 => x"8b168480",
   866 => x"8080af2d",
   867 => x"98065877",
   868 => x"8187388b",
   869 => x"537c5275",
   870 => x"51848080",
   871 => x"8fd02d83",
   872 => x"ffe08008",
   873 => x"80f3389c",
   874 => x"16085184",
   875 => x"80808cb1",
   876 => x"2d83ffe0",
   877 => x"8008841c",
   878 => x"0c9a1684",
   879 => x"8080809a",
   880 => x"2d518480",
   881 => x"808ce32d",
   882 => x"83ffe080",
   883 => x"0883ffe0",
   884 => x"80085555",
   885 => x"83fff5e0",
   886 => x"08802ea0",
   887 => x"38941684",
   888 => x"8080809a",
   889 => x"2d518480",
   890 => x"808ce32d",
   891 => x"83ffe080",
   892 => x"08902b83",
   893 => x"fff00a06",
   894 => x"70165154",
   895 => x"73881c0c",
   896 => x"777b0c7c",
   897 => x"52848080",
   898 => x"a4885184",
   899 => x"80808184",
   900 => x"2d7b5484",
   901 => x"80809cf4",
   902 => x"04811a5a",
   903 => x"8480809a",
   904 => x"ad0483ff",
   905 => x"f5e00880",
   906 => x"2e80c738",
   907 => x"76518480",
   908 => x"8098cc2d",
   909 => x"83ffe080",
   910 => x"0883ffe0",
   911 => x"80085384",
   912 => x"8080a49c",
   913 => x"52578480",
   914 => x"8081842d",
   915 => x"7680ffff",
   916 => x"fff80654",
   917 => x"7380ffff",
   918 => x"fff82e96",
   919 => x"38fe1783",
   920 => x"fff5e808",
   921 => x"2983fff5",
   922 => x"f0080555",
   923 => x"8480809a",
   924 => x"ab048054",
   925 => x"7383ffe0",
   926 => x"800c02b4",
   927 => x"050d0402",
   928 => x"e4050d78",
   929 => x"7a715483",
   930 => x"fff5bc53",
   931 => x"55558480",
   932 => x"8099ef2d",
   933 => x"83ffe080",
   934 => x"0881ff06",
   935 => x"5372802e",
   936 => x"81883884",
   937 => x"8080a4b4",
   938 => x"51848080",
   939 => x"84922d83",
   940 => x"fff5c008",
   941 => x"83ff0589",
   942 => x"2a578070",
   943 => x"56567577",
   944 => x"25818738",
   945 => x"83fff5c4",
   946 => x"08fe0583",
   947 => x"fff5e808",
   948 => x"2983fff5",
   949 => x"f0081176",
   950 => x"83fff5dc",
   951 => x"08060575",
   952 => x"54525384",
   953 => x"80808afd",
   954 => x"2d83ffe0",
   955 => x"8008802e",
   956 => x"80cc3881",
   957 => x"157083ff",
   958 => x"f5dc0806",
   959 => x"54557297",
   960 => x"3883fff5",
   961 => x"c4085184",
   962 => x"808098cc",
   963 => x"2d83ffe0",
   964 => x"800883ff",
   965 => x"f5c40c84",
   966 => x"80148117",
   967 => x"57547676",
   968 => x"24ffa138",
   969 => x"8480809e",
   970 => x"ca047452",
   971 => x"848080a4",
   972 => x"d0518480",
   973 => x"8081842d",
   974 => x"8480809e",
   975 => x"cc0483ff",
   976 => x"e0800853",
   977 => x"8480809e",
   978 => x"cc048153",
   979 => x"7283ffe0",
   980 => x"800c029c",
   981 => x"050d0483",
   982 => x"ffe08c08",
   983 => x"0283ffe0",
   984 => x"8c0cff3d",
   985 => x"0d800b83",
   986 => x"ffe08c08",
   987 => x"fc050c83",
   988 => x"ffe08c08",
   989 => x"88050881",
   990 => x"06ff1170",
   991 => x"097083ff",
   992 => x"e08c088c",
   993 => x"05080683",
   994 => x"ffe08c08",
   995 => x"fc050811",
   996 => x"83ffe08c",
   997 => x"08fc050c",
   998 => x"83ffe08c",
   999 => x"08880508",
  1000 => x"812a83ff",
  1001 => x"e08c0888",
  1002 => x"050c83ff",
  1003 => x"e08c088c",
  1004 => x"05081083",
  1005 => x"ffe08c08",
  1006 => x"8c050c51",
  1007 => x"51515183",
  1008 => x"ffe08c08",
  1009 => x"88050880",
  1010 => x"2e8438ff",
  1011 => x"a23983ff",
  1012 => x"e08c08fc",
  1013 => x"05087083",
  1014 => x"ffe0800c",
  1015 => x"51833d0d",
  1016 => x"83ffe08c",
  1017 => x"0c040000",
  1018 => x"00ffffff",
  1019 => x"ff00ffff",
  1020 => x"ffff00ff",
  1021 => x"ffffff00",
  1022 => x"436d645f",
  1023 => x"696e6974",
  1024 => x"0a000000",
  1025 => x"636d645f",
  1026 => x"434d4438",
  1027 => x"20726573",
  1028 => x"706f6e73",
  1029 => x"653a2025",
  1030 => x"640a0000",
  1031 => x"53444843",
  1032 => x"20496e69",
  1033 => x"7469616c",
  1034 => x"697a6174",
  1035 => x"696f6e20",
  1036 => x"6572726f",
  1037 => x"72210a00",
  1038 => x"434d4438",
  1039 => x"5f342072",
  1040 => x"6573706f",
  1041 => x"6e73653a",
  1042 => x"2025640a",
  1043 => x"00000000",
  1044 => x"434d4435",
  1045 => x"38202564",
  1046 => x"0a202000",
  1047 => x"434d4435",
  1048 => x"385f3220",
  1049 => x"25640a20",
  1050 => x"20000000",
  1051 => x"52656164",
  1052 => x"20636f6d",
  1053 => x"6d616e64",
  1054 => x"20666169",
  1055 => x"6c656420",
  1056 => x"61742025",
  1057 => x"64202825",
  1058 => x"64290a00",
  1059 => x"496e6974",
  1060 => x"69616c69",
  1061 => x"7a696e67",
  1062 => x"20534420",
  1063 => x"63617264",
  1064 => x"0a000000",
  1065 => x"48756e74",
  1066 => x"696e6720",
  1067 => x"666f7220",
  1068 => x"70617274",
  1069 => x"6974696f",
  1070 => x"6e0a0000",
  1071 => x"4d414e49",
  1072 => x"46455354",
  1073 => x"4d535400",
  1074 => x"50617273",
  1075 => x"696e6720",
  1076 => x"6d616e69",
  1077 => x"66657374",
  1078 => x"0a000000",
  1079 => x"52657475",
  1080 => x"726e696e",
  1081 => x"670a0000",
  1082 => x"52656164",
  1083 => x"696e6720",
  1084 => x"4d42520a",
  1085 => x"00000000",
  1086 => x"52656164",
  1087 => x"206f6620",
  1088 => x"4d425220",
  1089 => x"6661696c",
  1090 => x"65640a00",
  1091 => x"4d425220",
  1092 => x"73756363",
  1093 => x"65737366",
  1094 => x"756c6c79",
  1095 => x"20726561",
  1096 => x"640a0000",
  1097 => x"46415431",
  1098 => x"36202020",
  1099 => x"00000000",
  1100 => x"46415433",
  1101 => x"32202020",
  1102 => x"00000000",
  1103 => x"50617274",
  1104 => x"6974696f",
  1105 => x"6e636f75",
  1106 => x"6e742025",
  1107 => x"640a0000",
  1108 => x"4e6f2070",
  1109 => x"61727469",
  1110 => x"74696f6e",
  1111 => x"20736967",
  1112 => x"6e617475",
  1113 => x"72652066",
  1114 => x"6f756e64",
  1115 => x"0a000000",
  1116 => x"52656164",
  1117 => x"696e6720",
  1118 => x"626f6f74",
  1119 => x"20736563",
  1120 => x"746f7220",
  1121 => x"25640a00",
  1122 => x"52656164",
  1123 => x"20626f6f",
  1124 => x"74207365",
  1125 => x"63746f72",
  1126 => x"2066726f",
  1127 => x"6d206669",
  1128 => x"72737420",
  1129 => x"70617274",
  1130 => x"6974696f",
  1131 => x"6e0a0000",
  1132 => x"48756e74",
  1133 => x"696e6720",
  1134 => x"666f7220",
  1135 => x"66696c65",
  1136 => x"73797374",
  1137 => x"656d0a00",
  1138 => x"556e7375",
  1139 => x"70706f72",
  1140 => x"74656420",
  1141 => x"70617274",
  1142 => x"6974696f",
  1143 => x"6e207479",
  1144 => x"7065210d",
  1145 => x"00000000",
  1146 => x"52656164",
  1147 => x"696e6720",
  1148 => x"64697265",
  1149 => x"63746f72",
  1150 => x"79207365",
  1151 => x"63746f72",
  1152 => x"2025640a",
  1153 => x"00000000",
  1154 => x"66696c65",
  1155 => x"20222573",
  1156 => x"2220666f",
  1157 => x"756e640d",
  1158 => x"00000000",
  1159 => x"47657446",
  1160 => x"41544c69",
  1161 => x"6e6b2072",
  1162 => x"65747572",
  1163 => x"6e656420",
  1164 => x"25640a00",
  1165 => x"4f70656e",
  1166 => x"65642066",
  1167 => x"696c652c",
  1168 => x"206c6f61",
  1169 => x"64696e67",
  1170 => x"2e2e2e0a",
  1171 => x"00000000",
  1172 => x"43616e27",
  1173 => x"74206f70",
  1174 => x"656e2025",
  1175 => x"730a0000",
	others => x"00000000"
);

begin

process (clk)
begin
	if (clk'event and clk = '1') then
		if (from_zpu.memAWriteEnable = '1') and (from_zpu.memBWriteEnable = '1') and (from_zpu.memAAddr=from_zpu.memBAddr) and (from_zpu.memAWrite/=from_zpu.memBWrite) then
			report "write collision" severity failure;
		end if;
	
		if (from_zpu.memAWriteEnable = '1') then
			ram(to_integer(unsigned(from_zpu.memAAddr(maxAddrBitBRAM downto 2)))) := from_zpu.memAWrite;
			to_zpu.memARead <= from_zpu.memAWrite;
		else
			to_zpu.memARead <= ram(to_integer(unsigned(from_zpu.memAAddr(maxAddrBitBRAM downto 2))));
		end if;
	end if;
end process;

process (clk)
begin
	if (clk'event and clk = '1') then
		if (from_zpu.memBWriteEnable = '1') then
			ram(to_integer(unsigned(from_zpu.memBAddr(maxAddrBitBRAM downto 2)))) := from_zpu.memBWrite;
			to_zpu.memBRead <= from_zpu.memBWrite;
		else
			to_zpu.memBRead <= ram(to_integer(unsigned(from_zpu.memBAddr(maxAddrBitBRAM downto 2))));
		end if;
	end if;
end process;


end arch;

