-- ZPU
--
-- Copyright 2004-2008 oharboe - �yvind Harboe - oyvind.harboe@zylin.com
-- Modified by Alastair M. Robinson for the ZPUFlex project.
--
-- The FreeBSD license
-- 
-- Redistribution and use in source and binary forms, with or without
-- modification, are permitted provided that the following conditions
-- are met:
-- 
-- 1. Redistributions of source code must retain the above copyright
--    notice, this list of conditions and the following disclaimer.
-- 2. Redistributions in binary form must reproduce the above
--    copyright notice, this list of conditions and the following
--    disclaimer in the documentation and/or other materials
--    provided with the distribution.
-- 
-- THIS SOFTWARE IS PROVIDED BY THE ZPU PROJECT ``AS IS'' AND ANY
-- EXPRESS OR IMPLIED WARRANTIES, INCLUDING, BUT NOT LIMITED TO,
-- THE IMPLIED WARRANTIES OF MERCHANTABILITY AND FITNESS FOR A
-- PARTICULAR PURPOSE ARE DISCLAIMED. IN NO EVENT SHALL THE
-- ZPU PROJECT OR CONTRIBUTORS BE LIABLE FOR ANY DIRECT,
-- INDIRECT, INCIDENTAL, SPECIAL, EXEMPLARY, OR CONSEQUENTIAL DAMAGES
-- (INCLUDING, BUT NOT LIMITED TO, PROCUREMENT OF SUBSTITUTE GOODS
-- OR SERVICES; LOSS OF USE, DATA, OR PROFITS; OR BUSINESS INTERRUPTION)
-- HOWEVER CAUSED AND ON ANY THEORY OF LIABILITY, WHETHER IN CONTRACT,
-- STRICT LIABILITY, OR TORT (INCLUDING NEGLIGENCE OR OTHERWISE)
-- ARISING IN ANY WAY OUT OF THE USE OF THIS SOFTWARE, EVEN IF
-- ADVISED OF THE POSSIBILITY OF SUCH DAMAGE.
-- 
-- The views and conclusions contained in the software and documentation
-- are those of the authors and should not be interpreted as representing
-- official policies, either expressed or implied, of the ZPU Project.

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;


library work;
use work.zpu_config.all;
use work.zpupkg.all;

entity SDRAMTest_ROM is
generic
	(
		maxAddrBitBRAM : integer := maxAddrBitBRAMLimit -- Specify your actual ROM size to save LEs and unnecessary block RAM usage.
	);
port (
	clk : in std_logic;
	areset : in std_logic := '0';
	from_zpu : in ZPU_ToROM;
	to_zpu : out ZPU_FromROM
);
end SDRAMTest_ROM;

architecture arch of SDRAMTest_ROM is

type ram_type is array(natural range 0 to ((2**(maxAddrBitBRAM+1))/4)-1) of std_logic_vector(wordSize-1 downto 0);

shared variable ram : ram_type :=
(
     0 => x"84808080",
     1 => x"ed040000",
     2 => x"00000000",
     3 => x"84808080",
     4 => x"880d8004",
     5 => x"84808080",
     6 => x"940471fd",
     7 => x"06087283",
     8 => x"06098105",
     9 => x"8205832b",
    10 => x"2a83ffff",
    11 => x"06520471",
    12 => x"fc060872",
    13 => x"83060981",
    14 => x"05830510",
    15 => x"10102a81",
    16 => x"ff065204",
    17 => x"71fc0608",
    18 => x"8480808f",
    19 => x"f4738306",
    20 => x"10100508",
    21 => x"067381ff",
    22 => x"06738306",
    23 => x"09810583",
    24 => x"05101010",
    25 => x"2b0772fc",
    26 => x"060c5151",
    27 => x"04028405",
    28 => x"84808080",
    29 => x"880c8480",
    30 => x"8080940b",
    31 => x"8480808c",
    32 => x"e1040000",
    33 => x"02c0050d",
    34 => x"0280c405",
    35 => x"84808096",
    36 => x"e05c5c80",
    37 => x"7c708405",
    38 => x"5e08715f",
    39 => x"5f587d70",
    40 => x"84055f08",
    41 => x"57805976",
    42 => x"982a7788",
    43 => x"2b585574",
    44 => x"802e82a9",
    45 => x"387c802e",
    46 => x"80c53880",
    47 => x"5d7480e4",
    48 => x"2e81bb38",
    49 => x"7480e426",
    50 => x"80f13874",
    51 => x"80e32e80",
    52 => x"c838a551",
    53 => x"84808084",
    54 => x"912d7451",
    55 => x"84808084",
    56 => x"912d8218",
    57 => x"58811959",
    58 => x"837925ff",
    59 => x"ba3874ff",
    60 => x"ad387e84",
    61 => x"80809680",
    62 => x"0c0280c0",
    63 => x"050d0474",
    64 => x"a52e0981",
    65 => x"069b3881",
    66 => x"0b811a5a",
    67 => x"5d837925",
    68 => x"ff953884",
    69 => x"808081ee",
    70 => x"047b841d",
    71 => x"7108575d",
    72 => x"54745184",
    73 => x"80808491",
    74 => x"2d811881",
    75 => x"1a5a5883",
    76 => x"7925fef3",
    77 => x"38848080",
    78 => x"81ee0474",
    79 => x"80f32e09",
    80 => x"8106ff8e",
    81 => x"387b841d",
    82 => x"71087054",
    83 => x"5d5d5384",
    84 => x"808084b6",
    85 => x"2d800bff",
    86 => x"11545280",
    87 => x"7225ff85",
    88 => x"387a7081",
    89 => x"055c3370",
    90 => x"52558480",
    91 => x"8084912d",
    92 => x"811873ff",
    93 => x"15555358",
    94 => x"84808082",
    95 => x"db047b84",
    96 => x"1d71087f",
    97 => x"5d555d52",
    98 => x"80732480",
    99 => x"f1387280",
   100 => x"2e80d738",
   101 => x"8756729c",
   102 => x"2a73842b",
   103 => x"54527180",
   104 => x"2e833881",
   105 => x"5ab71254",
   106 => x"71892484",
   107 => x"38b01254",
   108 => x"799538ff",
   109 => x"16567580",
   110 => x"25dc3880",
   111 => x"0bff1154",
   112 => x"52848080",
   113 => x"82db0473",
   114 => x"51848080",
   115 => x"84912dff",
   116 => x"16567580",
   117 => x"25c03884",
   118 => x"808083bb",
   119 => x"04778480",
   120 => x"8096800c",
   121 => x"0280c005",
   122 => x"0d04b051",
   123 => x"84808084",
   124 => x"912d800b",
   125 => x"ff115452",
   126 => x"84808082",
   127 => x"db04ad51",
   128 => x"84808084",
   129 => x"912d7209",
   130 => x"81055384",
   131 => x"8080838e",
   132 => x"0402f805",
   133 => x"0d7352c0",
   134 => x"0870882a",
   135 => x"70810651",
   136 => x"51517080",
   137 => x"2ef13871",
   138 => x"c00c7184",
   139 => x"80809680",
   140 => x"0c028805",
   141 => x"0d0402e8",
   142 => x"050d8078",
   143 => x"57557570",
   144 => x"84055708",
   145 => x"53805472",
   146 => x"982a7388",
   147 => x"2b545271",
   148 => x"802ea238",
   149 => x"c0087088",
   150 => x"2a708106",
   151 => x"51515170",
   152 => x"802ef138",
   153 => x"71c00c81",
   154 => x"15811555",
   155 => x"55837425",
   156 => x"d63871ca",
   157 => x"38748480",
   158 => x"8096800c",
   159 => x"0298050d",
   160 => x"0402f405",
   161 => x"0d747652",
   162 => x"53807125",
   163 => x"90387052",
   164 => x"72708405",
   165 => x"5408ff13",
   166 => x"535171f4",
   167 => x"38028c05",
   168 => x"0d0402d4",
   169 => x"050d7c7e",
   170 => x"5c58810b",
   171 => x"84808090",
   172 => x"84585a83",
   173 => x"59760878",
   174 => x"0c770877",
   175 => x"08565473",
   176 => x"752e9438",
   177 => x"77085374",
   178 => x"52848080",
   179 => x"90945184",
   180 => x"80808184",
   181 => x"2d805a77",
   182 => x"56807b25",
   183 => x"90387a55",
   184 => x"75708405",
   185 => x"5708ff16",
   186 => x"565474f4",
   187 => x"38770877",
   188 => x"08565675",
   189 => x"752e9438",
   190 => x"77085374",
   191 => x"52848080",
   192 => x"90d45184",
   193 => x"80808184",
   194 => x"2d805aff",
   195 => x"19841858",
   196 => x"59788025",
   197 => x"ff9f3879",
   198 => x"84808096",
   199 => x"800c02ac",
   200 => x"050d0402",
   201 => x"e4050d78",
   202 => x"7a555681",
   203 => x"5785aad5",
   204 => x"aad5760c",
   205 => x"fad5aad5",
   206 => x"aa0b8c17",
   207 => x"0ccc7634",
   208 => x"b30b8f17",
   209 => x"34750853",
   210 => x"72fce2d5",
   211 => x"aad52e92",
   212 => x"38750852",
   213 => x"84808091",
   214 => x"94518480",
   215 => x"8081842d",
   216 => x"80578c16",
   217 => x"085574fa",
   218 => x"d5aad4b3",
   219 => x"2e93388c",
   220 => x"16085284",
   221 => x"808091d0",
   222 => x"51848080",
   223 => x"81842d80",
   224 => x"57755580",
   225 => x"74258e38",
   226 => x"74708405",
   227 => x"5608ff15",
   228 => x"555373f4",
   229 => x"38750854",
   230 => x"73fce2d5",
   231 => x"aad52e92",
   232 => x"38750852",
   233 => x"84808092",
   234 => x"8c518480",
   235 => x"8081842d",
   236 => x"80578c16",
   237 => x"085372fa",
   238 => x"d5aad4b3",
   239 => x"2e93388c",
   240 => x"16085284",
   241 => x"808092c8",
   242 => x"51848080",
   243 => x"81842d80",
   244 => x"57768480",
   245 => x"8096800c",
   246 => x"029c050d",
   247 => x"0402c405",
   248 => x"0d605b80",
   249 => x"62908080",
   250 => x"29ff0584",
   251 => x"80809384",
   252 => x"53405a84",
   253 => x"80808184",
   254 => x"2d80e1b3",
   255 => x"5780fe5e",
   256 => x"ae518480",
   257 => x"8084912d",
   258 => x"76107096",
   259 => x"2a810656",
   260 => x"5774802e",
   261 => x"85387681",
   262 => x"07577695",
   263 => x"2a810658",
   264 => x"77802e85",
   265 => x"38768132",
   266 => x"57787707",
   267 => x"7f06775e",
   268 => x"598fffff",
   269 => x"5876bfff",
   270 => x"ff06707a",
   271 => x"32822b7c",
   272 => x"11515776",
   273 => x"0c761070",
   274 => x"962a8106",
   275 => x"56577480",
   276 => x"2e853876",
   277 => x"81075776",
   278 => x"952a8106",
   279 => x"5574802e",
   280 => x"85387681",
   281 => x"3257ff18",
   282 => x"58778025",
   283 => x"c8387c57",
   284 => x"8fffff58",
   285 => x"76bfffff",
   286 => x"06707a32",
   287 => x"822b7c05",
   288 => x"7008575e",
   289 => x"5674762e",
   290 => x"80ea3880",
   291 => x"7a538480",
   292 => x"80939452",
   293 => x"5c848080",
   294 => x"81842d74",
   295 => x"54755375",
   296 => x"52848080",
   297 => x"93a85184",
   298 => x"80808184",
   299 => x"2d7b5a76",
   300 => x"1070962a",
   301 => x"81065757",
   302 => x"75802e85",
   303 => x"38768107",
   304 => x"5776952a",
   305 => x"81065574",
   306 => x"802e8538",
   307 => x"76813257",
   308 => x"ff185877",
   309 => x"8025ff9c",
   310 => x"38ff1e5e",
   311 => x"7dfea138",
   312 => x"8a518480",
   313 => x"8084912d",
   314 => x"7b848080",
   315 => x"96800c02",
   316 => x"bc050d04",
   317 => x"811a5a84",
   318 => x"808089af",
   319 => x"0402cc05",
   320 => x"0d7e605e",
   321 => x"58815a80",
   322 => x"5b80c07a",
   323 => x"585c85ad",
   324 => x"a989bb78",
   325 => x"0c795981",
   326 => x"56975576",
   327 => x"7607822b",
   328 => x"78115154",
   329 => x"85ada989",
   330 => x"bb740c75",
   331 => x"10ff1656",
   332 => x"56748025",
   333 => x"e6387610",
   334 => x"811a5a57",
   335 => x"987925d7",
   336 => x"38775680",
   337 => x"7d259038",
   338 => x"7c557570",
   339 => x"84055708",
   340 => x"ff165654",
   341 => x"74f43881",
   342 => x"57ff8787",
   343 => x"a5c3780c",
   344 => x"97597682",
   345 => x"2b781170",
   346 => x"085f5656",
   347 => x"7cff8787",
   348 => x"a5c32e80",
   349 => x"cc387408",
   350 => x"547385ad",
   351 => x"a989bb2e",
   352 => x"94388075",
   353 => x"08547653",
   354 => x"84808093",
   355 => x"d0525a84",
   356 => x"80808184",
   357 => x"2d7610ff",
   358 => x"1a5a5778",
   359 => x"8025c338",
   360 => x"7a822b56",
   361 => x"75b1387b",
   362 => x"52848080",
   363 => x"93f05184",
   364 => x"80808184",
   365 => x"2d7b8480",
   366 => x"8096800c",
   367 => x"02b4050d",
   368 => x"047a7707",
   369 => x"7710ff1b",
   370 => x"5b585b78",
   371 => x"8025ff92",
   372 => x"38848080",
   373 => x"8ba00475",
   374 => x"52848080",
   375 => x"94ac5184",
   376 => x"80808184",
   377 => x"2d75992a",
   378 => x"81328106",
   379 => x"70098105",
   380 => x"71077009",
   381 => x"709f2c7d",
   382 => x"0679109f",
   383 => x"fffffc06",
   384 => x"60812a41",
   385 => x"5a5d5758",
   386 => x"5975da38",
   387 => x"79098105",
   388 => x"707b079f",
   389 => x"2a55567b",
   390 => x"bf268438",
   391 => x"739d3881",
   392 => x"70538480",
   393 => x"8093f052",
   394 => x"5c848080",
   395 => x"81842d7b",
   396 => x"84808096",
   397 => x"800c02b4",
   398 => x"050d0484",
   399 => x"808094c4",
   400 => x"51848080",
   401 => x"81842d7b",
   402 => x"52848080",
   403 => x"93f05184",
   404 => x"80808184",
   405 => x"2d7b8480",
   406 => x"8096800c",
   407 => x"02b4050d",
   408 => x"0402dc05",
   409 => x"0d810b84",
   410 => x"80809084",
   411 => x"58588359",
   412 => x"7608800c",
   413 => x"80087708",
   414 => x"56547375",
   415 => x"2e943880",
   416 => x"08537452",
   417 => x"84808090",
   418 => x"94518480",
   419 => x"8081842d",
   420 => x"80588070",
   421 => x"57557570",
   422 => x"84055708",
   423 => x"81165654",
   424 => x"a0807524",
   425 => x"f1388008",
   426 => x"77085656",
   427 => x"75752e94",
   428 => x"38800853",
   429 => x"74528480",
   430 => x"8090d451",
   431 => x"84808081",
   432 => x"842d8058",
   433 => x"ff198418",
   434 => x"58597880",
   435 => x"25ffa138",
   436 => x"77802e8d",
   437 => x"38848080",
   438 => x"95905184",
   439 => x"80808184",
   440 => x"2d815785",
   441 => x"aad5aad5",
   442 => x"0b800cfa",
   443 => x"d5aad5aa",
   444 => x"0b8c0ccc",
   445 => x"0b8034b3",
   446 => x"0b8f3480",
   447 => x"085574fc",
   448 => x"e2d5aad5",
   449 => x"2e923880",
   450 => x"08528480",
   451 => x"80919451",
   452 => x"84808081",
   453 => x"842d8057",
   454 => x"8c085877",
   455 => x"fad5aad4",
   456 => x"b32e9238",
   457 => x"8c085284",
   458 => x"808091d0",
   459 => x"51848080",
   460 => x"81842d80",
   461 => x"57807057",
   462 => x"55757084",
   463 => x"05570881",
   464 => x"165654a0",
   465 => x"807524f1",
   466 => x"38800859",
   467 => x"78fce2d5",
   468 => x"aad52e92",
   469 => x"38800852",
   470 => x"84808092",
   471 => x"8c518480",
   472 => x"8081842d",
   473 => x"80578c08",
   474 => x"5473fad5",
   475 => x"aad4b32e",
   476 => x"80ea388c",
   477 => x"08528480",
   478 => x"8092c851",
   479 => x"84808081",
   480 => x"842da080",
   481 => x"52805184",
   482 => x"808089fd",
   483 => x"2d848080",
   484 => x"96800854",
   485 => x"84808096",
   486 => x"8008802e",
   487 => x"8d388480",
   488 => x"8095b451",
   489 => x"84808081",
   490 => x"842d7352",
   491 => x"80518480",
   492 => x"8087dd2d",
   493 => x"84808096",
   494 => x"8008802e",
   495 => x"fda73884",
   496 => x"808095cc",
   497 => x"51848080",
   498 => x"81842d81",
   499 => x"0b848080",
   500 => x"90845858",
   501 => x"83598480",
   502 => x"808cf004",
   503 => x"76802eff",
   504 => x"a1388480",
   505 => x"8095e451",
   506 => x"84808081",
   507 => x"842d8480",
   508 => x"808f8204",
   509 => x"00ffffff",
   510 => x"ff00ffff",
   511 => x"ffff00ff",
   512 => x"ffffff00",
   513 => x"00000000",
   514 => x"55555555",
   515 => x"aaaaaaaa",
   516 => x"ffffffff",
   517 => x"53616e69",
   518 => x"74792063",
   519 => x"6865636b",
   520 => x"20666169",
   521 => x"6c656420",
   522 => x"28626566",
   523 => x"6f726520",
   524 => x"63616368",
   525 => x"65207265",
   526 => x"66726573",
   527 => x"6829206f",
   528 => x"6e203078",
   529 => x"25642028",
   530 => x"676f7420",
   531 => x"30782564",
   532 => x"290a0000",
   533 => x"53616e69",
   534 => x"74792063",
   535 => x"6865636b",
   536 => x"20666169",
   537 => x"6c656420",
   538 => x"28616674",
   539 => x"65722063",
   540 => x"61636865",
   541 => x"20726566",
   542 => x"72657368",
   543 => x"29206f6e",
   544 => x"20307825",
   545 => x"64202867",
   546 => x"6f742030",
   547 => x"78256429",
   548 => x"0a000000",
   549 => x"42797465",
   550 => x"20636865",
   551 => x"636b2066",
   552 => x"61696c65",
   553 => x"64202862",
   554 => x"65666f72",
   555 => x"65206361",
   556 => x"63686520",
   557 => x"72656672",
   558 => x"65736829",
   559 => x"20617420",
   560 => x"30202867",
   561 => x"6f742030",
   562 => x"78256429",
   563 => x"0a000000",
   564 => x"42797465",
   565 => x"20636865",
   566 => x"636b2066",
   567 => x"61696c65",
   568 => x"64202862",
   569 => x"65666f72",
   570 => x"65206361",
   571 => x"63686520",
   572 => x"72656672",
   573 => x"65736829",
   574 => x"20617420",
   575 => x"33202867",
   576 => x"6f742030",
   577 => x"78256429",
   578 => x"0a000000",
   579 => x"42797465",
   580 => x"20636865",
   581 => x"636b2066",
   582 => x"61696c65",
   583 => x"64202861",
   584 => x"66746572",
   585 => x"20636163",
   586 => x"68652072",
   587 => x"65667265",
   588 => x"73682920",
   589 => x"61742030",
   590 => x"2028676f",
   591 => x"74203078",
   592 => x"2564290a",
   593 => x"00000000",
   594 => x"42797465",
   595 => x"20636865",
   596 => x"636b2066",
   597 => x"61696c65",
   598 => x"64202861",
   599 => x"66746572",
   600 => x"20636163",
   601 => x"68652072",
   602 => x"65667265",
   603 => x"73682920",
   604 => x"61742033",
   605 => x"2028676f",
   606 => x"74203078",
   607 => x"2564290a",
   608 => x"00000000",
   609 => x"43686563",
   610 => x"6b696e67",
   611 => x"206d656d",
   612 => x"6f727900",
   613 => x"30782564",
   614 => x"20676f6f",
   615 => x"64207265",
   616 => x"6164732c",
   617 => x"20000000",
   618 => x"4572726f",
   619 => x"72206174",
   620 => x"20307825",
   621 => x"642c2065",
   622 => x"78706563",
   623 => x"74656420",
   624 => x"30782564",
   625 => x"2c20676f",
   626 => x"74203078",
   627 => x"25640a00",
   628 => x"42616420",
   629 => x"64617461",
   630 => x"20666f75",
   631 => x"6e642061",
   632 => x"74203078",
   633 => x"25642028",
   634 => x"30782564",
   635 => x"290a0000",
   636 => x"53445241",
   637 => x"4d207369",
   638 => x"7a652028",
   639 => x"61737375",
   640 => x"6d696e67",
   641 => x"206e6f20",
   642 => x"61646472",
   643 => x"65737320",
   644 => x"6661756c",
   645 => x"74732920",
   646 => x"69732030",
   647 => x"78256420",
   648 => x"6d656761",
   649 => x"62797465",
   650 => x"730a0000",
   651 => x"416c6961",
   652 => x"73657320",
   653 => x"666f756e",
   654 => x"64206174",
   655 => x"20307825",
   656 => x"640a0000",
   657 => x"28416c69",
   658 => x"61736573",
   659 => x"2070726f",
   660 => x"6261626c",
   661 => x"79207369",
   662 => x"6d706c79",
   663 => x"20696e64",
   664 => x"69636174",
   665 => x"65207468",
   666 => x"61742052",
   667 => x"414d0a69",
   668 => x"7320736d",
   669 => x"616c6c65",
   670 => x"72207468",
   671 => x"616e2036",
   672 => x"34206d65",
   673 => x"67616279",
   674 => x"74657329",
   675 => x"0a000000",
   676 => x"46697273",
   677 => x"74207374",
   678 => x"61676520",
   679 => x"73616e69",
   680 => x"74792063",
   681 => x"6865636b",
   682 => x"20706173",
   683 => x"7365642e",
   684 => x"0a000000",
   685 => x"41646472",
   686 => x"65737320",
   687 => x"63686563",
   688 => x"6b207061",
   689 => x"73736564",
   690 => x"2e0a0000",
   691 => x"4c465352",
   692 => x"20636865",
   693 => x"636b2070",
   694 => x"61737365",
   695 => x"642e0a0a",
   696 => x"00000000",
   697 => x"42797465",
   698 => x"20286471",
   699 => x"6d292063",
   700 => x"6865636b",
   701 => x"20706173",
   702 => x"7365640a",
   703 => x"00000000",
	others => x"00000000"
);

begin

process (clk)
begin
	if (clk'event and clk = '1') then
		if (from_zpu.memAWriteEnable = '1') and (from_zpu.memBWriteEnable = '1') and (from_zpu.memAAddr=from_zpu.memBAddr) and (from_zpu.memAWrite/=from_zpu.memBWrite) then
			report "write collision" severity failure;
		end if;
	
		if (from_zpu.memAWriteEnable = '1') then
			ram(to_integer(unsigned(from_zpu.memAAddr(maxAddrBitBRAM downto 2)))) := from_zpu.memAWrite;
			to_zpu.memARead <= from_zpu.memAWrite;
		else
			to_zpu.memARead <= ram(to_integer(unsigned(from_zpu.memAAddr(maxAddrBitBRAM downto 2))));
		end if;
	end if;
end process;

process (clk)
begin
	if (clk'event and clk = '1') then
		if (from_zpu.memBWriteEnable = '1') then
			ram(to_integer(unsigned(from_zpu.memBAddr(maxAddrBitBRAM downto 2)))) := from_zpu.memBWrite;
			to_zpu.memBRead <= from_zpu.memBWrite;
		else
			to_zpu.memBRead <= ram(to_integer(unsigned(from_zpu.memBAddr(maxAddrBitBRAM downto 2))));
		end if;
	end if;
end process;


end arch;

