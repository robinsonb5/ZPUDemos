-- ZPU
--
-- Copyright 2004-2008 oharboe - �yvind Harboe - oyvind.harboe@zylin.com
-- Modified by Alastair M. Robinson for the ZPUFlex project.
--
-- The FreeBSD license
-- 
-- Redistribution and use in source and binary forms, with or without
-- modification, are permitted provided that the following conditions
-- are met:
-- 
-- 1. Redistributions of source code must retain the above copyright
--    notice, this list of conditions and the following disclaimer.
-- 2. Redistributions in binary form must reproduce the above
--    copyright notice, this list of conditions and the following
--    disclaimer in the documentation and/or other materials
--    provided with the distribution.
-- 
-- THIS SOFTWARE IS PROVIDED BY THE ZPU PROJECT ``AS IS'' AND ANY
-- EXPRESS OR IMPLIED WARRANTIES, INCLUDING, BUT NOT LIMITED TO,
-- THE IMPLIED WARRANTIES OF MERCHANTABILITY AND FITNESS FOR A
-- PARTICULAR PURPOSE ARE DISCLAIMED. IN NO EVENT SHALL THE
-- ZPU PROJECT OR CONTRIBUTORS BE LIABLE FOR ANY DIRECT,
-- INDIRECT, INCIDENTAL, SPECIAL, EXEMPLARY, OR CONSEQUENTIAL DAMAGES
-- (INCLUDING, BUT NOT LIMITED TO, PROCUREMENT OF SUBSTITUTE GOODS
-- OR SERVICES; LOSS OF USE, DATA, OR PROFITS; OR BUSINESS INTERRUPTION)
-- HOWEVER CAUSED AND ON ANY THEORY OF LIABILITY, WHETHER IN CONTRACT,
-- STRICT LIABILITY, OR TORT (INCLUDING NEGLIGENCE OR OTHERWISE)
-- ARISING IN ANY WAY OUT OF THE USE OF THIS SOFTWARE, EVEN IF
-- ADVISED OF THE POSSIBILITY OF SUCH DAMAGE.
-- 
-- The views and conclusions contained in the software and documentation
-- are those of the authors and should not be interpreted as representing
-- official policies, either expressed or implied, of the ZPU Project.

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;


library work;
use work.zpupkg.all;

entity SDBootstrap_ROM is
generic
	(
		maxAddrBitBRAM : integer := maxAddrBitBRAMLimit -- Specify your actual ROM size to save LEs and unnecessary block RAM usage.
	);
port (
	clk : in std_logic;
	areset : in std_logic := '0';
	from_zpu : in ZPU_ToROM;
	to_zpu : out ZPU_FromROM
);
end SDBootstrap_ROM;

architecture arch of SDBootstrap_ROM is

type ram_type is array(natural range 0 to ((2**(maxAddrBitBRAM+1))/4)-1) of std_logic_vector(wordSize-1 downto 0);

shared variable ram : ram_type :=
(
     0 => x"84808080",
     1 => x"8c0b8480",
     2 => x"8081e004",
     3 => x"84808080",
     4 => x"8c04ff0d",
     5 => x"80040400",
     6 => x"40000016",
     7 => x"00000000",
     8 => x"0b83ffe0",
     9 => x"80080b83",
    10 => x"ffe08408",
    11 => x"0b83ffe0",
    12 => x"88088480",
    13 => x"80809808",
    14 => x"2d0b83ff",
    15 => x"e0880c0b",
    16 => x"83ffe084",
    17 => x"0c0b83ff",
    18 => x"e0800c04",
    19 => x"00000000",
    20 => x"00000000",
    21 => x"00000000",
    22 => x"00000000",
    23 => x"00000000",
    24 => x"71fd0608",
    25 => x"72830609",
    26 => x"81058205",
    27 => x"832b2a83",
    28 => x"ffff0652",
    29 => x"0471fc06",
    30 => x"08728306",
    31 => x"09810583",
    32 => x"05101010",
    33 => x"2a81ff06",
    34 => x"520471fd",
    35 => x"060883ff",
    36 => x"ff738306",
    37 => x"09810582",
    38 => x"05832b2b",
    39 => x"09067383",
    40 => x"ffff0673",
    41 => x"83060981",
    42 => x"05820583",
    43 => x"2b0b2b07",
    44 => x"72fc060c",
    45 => x"51510471",
    46 => x"fc060884",
    47 => x"8080a1d4",
    48 => x"73830610",
    49 => x"10050806",
    50 => x"7381ff06",
    51 => x"73830609",
    52 => x"81058305",
    53 => x"1010102b",
    54 => x"0772fc06",
    55 => x"0c515104",
    56 => x"83ffe080",
    57 => x"7083fff5",
    58 => x"f0278e38",
    59 => x"80717084",
    60 => x"05530c84",
    61 => x"808081e4",
    62 => x"04848080",
    63 => x"808c5184",
    64 => x"80808fd2",
    65 => x"0402ec05",
    66 => x"0d765380",
    67 => x"55727525",
    68 => x"8e38ad51",
    69 => x"84808085",
    70 => x"b32d7209",
    71 => x"81055372",
    72 => x"802ebe38",
    73 => x"8754729c",
    74 => x"2a73842b",
    75 => x"54527180",
    76 => x"2e833881",
    77 => x"55897225",
    78 => x"8a38b712",
    79 => x"52848080",
    80 => x"82c604b0",
    81 => x"12527480",
    82 => x"2e893871",
    83 => x"51848080",
    84 => x"85b32dff",
    85 => x"14547380",
    86 => x"25cc3884",
    87 => x"808082e9",
    88 => x"04b05184",
    89 => x"808085b3",
    90 => x"2d800b83",
    91 => x"ffe0800c",
    92 => x"0294050d",
    93 => x"0402c005",
    94 => x"0d0280c4",
    95 => x"05578070",
    96 => x"78708405",
    97 => x"5a087241",
    98 => x"5f5d587c",
    99 => x"7084055e",
   100 => x"085a805b",
   101 => x"79982a7a",
   102 => x"882b5b56",
   103 => x"75893877",
   104 => x"5f848080",
   105 => x"85a7047d",
   106 => x"802e81d3",
   107 => x"38805e75",
   108 => x"80e42e8a",
   109 => x"387580f8",
   110 => x"2e098106",
   111 => x"89387684",
   112 => x"1871085e",
   113 => x"58547580",
   114 => x"e42ea638",
   115 => x"7580e426",
   116 => x"8e387580",
   117 => x"e32e80d9",
   118 => x"38848080",
   119 => x"84bf0475",
   120 => x"80f32eb5",
   121 => x"387580f8",
   122 => x"2e8f3884",
   123 => x"808084bf",
   124 => x"048a5384",
   125 => x"808083fb",
   126 => x"04905383",
   127 => x"ffe0e052",
   128 => x"7b518480",
   129 => x"8082852d",
   130 => x"83ffe080",
   131 => x"0883ffe0",
   132 => x"e05a5584",
   133 => x"808084d8",
   134 => x"04768418",
   135 => x"71087054",
   136 => x"5b585484",
   137 => x"808085d7",
   138 => x"2d805584",
   139 => x"808084d8",
   140 => x"04768418",
   141 => x"71085858",
   142 => x"54848080",
   143 => x"858f04a5",
   144 => x"51848080",
   145 => x"85b32d75",
   146 => x"51848080",
   147 => x"85b32d82",
   148 => x"18588480",
   149 => x"80859a04",
   150 => x"74ff1656",
   151 => x"54807425",
   152 => x"b9387870",
   153 => x"81055a84",
   154 => x"808080f5",
   155 => x"2d705256",
   156 => x"84808085",
   157 => x"b32d8118",
   158 => x"58848080",
   159 => x"84d80475",
   160 => x"a52e0981",
   161 => x"06893881",
   162 => x"5e848080",
   163 => x"859a0475",
   164 => x"51848080",
   165 => x"85b32d81",
   166 => x"1858811b",
   167 => x"5b837b25",
   168 => x"fdf23875",
   169 => x"fde5387e",
   170 => x"83ffe080",
   171 => x"0c0280c0",
   172 => x"050d0402",
   173 => x"f8050d73",
   174 => x"52c00870",
   175 => x"882a7081",
   176 => x"06515151",
   177 => x"70802ef1",
   178 => x"3871c00c",
   179 => x"7183ffe0",
   180 => x"800c0288",
   181 => x"050d0402",
   182 => x"e8050d80",
   183 => x"78575575",
   184 => x"70840557",
   185 => x"08538054",
   186 => x"72982a73",
   187 => x"882b5452",
   188 => x"71802ea2",
   189 => x"38c00870",
   190 => x"882a7081",
   191 => x"06515151",
   192 => x"70802ef1",
   193 => x"3871c00c",
   194 => x"81158115",
   195 => x"55558374",
   196 => x"25d63871",
   197 => x"ca387483",
   198 => x"ffe0800c",
   199 => x"0298050d",
   200 => x"0402f405",
   201 => x"0dd45281",
   202 => x"ff720c71",
   203 => x"085381ff",
   204 => x"720c7288",
   205 => x"2b83fe80",
   206 => x"06720870",
   207 => x"81ff0651",
   208 => x"525381ff",
   209 => x"720c7271",
   210 => x"07882b72",
   211 => x"087081ff",
   212 => x"06515253",
   213 => x"81ff720c",
   214 => x"72710788",
   215 => x"2b720870",
   216 => x"81ff0672",
   217 => x"0783ffe0",
   218 => x"800c5253",
   219 => x"028c050d",
   220 => x"0402f405",
   221 => x"0d747671",
   222 => x"81ff06d4",
   223 => x"0c535383",
   224 => x"fff1a008",
   225 => x"85387189",
   226 => x"2b527198",
   227 => x"2ad40c71",
   228 => x"902a7081",
   229 => x"ff06d40c",
   230 => x"5171882a",
   231 => x"7081ff06",
   232 => x"d40c5171",
   233 => x"81ff06d4",
   234 => x"0c72902a",
   235 => x"7081ff06",
   236 => x"d40c51d4",
   237 => x"087081ff",
   238 => x"06515182",
   239 => x"b8bf5270",
   240 => x"81ff2e09",
   241 => x"81069438",
   242 => x"81ff0bd4",
   243 => x"0cd40870",
   244 => x"81ff06ff",
   245 => x"14545151",
   246 => x"71e53870",
   247 => x"83ffe080",
   248 => x"0c028c05",
   249 => x"0d0402fc",
   250 => x"050d81c7",
   251 => x"5181ff0b",
   252 => x"d40cff11",
   253 => x"51708025",
   254 => x"f4380284",
   255 => x"050d0402",
   256 => x"f0050d84",
   257 => x"808087e6",
   258 => x"2d819c9f",
   259 => x"53805287",
   260 => x"fc80f751",
   261 => x"84808086",
   262 => x"f12d83ff",
   263 => x"e0800854",
   264 => x"83ffe080",
   265 => x"08812e09",
   266 => x"8106ae38",
   267 => x"81ff0bd4",
   268 => x"0c820a52",
   269 => x"849c80e9",
   270 => x"51848080",
   271 => x"86f12d83",
   272 => x"ffe08008",
   273 => x"8e3881ff",
   274 => x"0bd40c73",
   275 => x"53848080",
   276 => x"88e00484",
   277 => x"808087e6",
   278 => x"2dff1353",
   279 => x"72ffae38",
   280 => x"7283ffe0",
   281 => x"800c0290",
   282 => x"050d0402",
   283 => x"f4050d81",
   284 => x"ff0bd40c",
   285 => x"848080a1",
   286 => x"e4518480",
   287 => x"8085d72d",
   288 => x"93538052",
   289 => x"87fc80c1",
   290 => x"51848080",
   291 => x"86f12d83",
   292 => x"ffe08008",
   293 => x"8e3881ff",
   294 => x"0bd40c81",
   295 => x"53848080",
   296 => x"89af0484",
   297 => x"808087e6",
   298 => x"2dff1353",
   299 => x"72d43872",
   300 => x"83ffe080",
   301 => x"0c028c05",
   302 => x"0d0402f0",
   303 => x"050d8480",
   304 => x"8087e62d",
   305 => x"83aa5284",
   306 => x"9c80c851",
   307 => x"84808086",
   308 => x"f12d83ff",
   309 => x"e0800883",
   310 => x"ffe08008",
   311 => x"53848080",
   312 => x"a1f05253",
   313 => x"84808082",
   314 => x"f52d7281",
   315 => x"2e098106",
   316 => x"a9388480",
   317 => x"8086a12d",
   318 => x"83ffe080",
   319 => x"0883ffff",
   320 => x"06537283",
   321 => x"aa2ebb38",
   322 => x"83ffe080",
   323 => x"08528480",
   324 => x"80a28851",
   325 => x"84808082",
   326 => x"f52d8480",
   327 => x"8088eb2d",
   328 => x"8480808a",
   329 => x"ba048154",
   330 => x"8480808b",
   331 => x"e5048480",
   332 => x"80a2a051",
   333 => x"84808082",
   334 => x"f52d8054",
   335 => x"8480808b",
   336 => x"e50481ff",
   337 => x"0bd40cb1",
   338 => x"53848080",
   339 => x"87ff2d83",
   340 => x"ffe08008",
   341 => x"802e80fe",
   342 => x"38805287",
   343 => x"fc80fa51",
   344 => x"84808086",
   345 => x"f12d83ff",
   346 => x"e0800880",
   347 => x"d73883ff",
   348 => x"e0800852",
   349 => x"848080a2",
   350 => x"bc518480",
   351 => x"8082f52d",
   352 => x"81ff0bd4",
   353 => x"0cd40870",
   354 => x"81ff0670",
   355 => x"54848080",
   356 => x"a2c85351",
   357 => x"53848080",
   358 => x"82f52d81",
   359 => x"ff0bd40c",
   360 => x"81ff0bd4",
   361 => x"0c81ff0b",
   362 => x"d40c81ff",
   363 => x"0bd40c72",
   364 => x"862a7081",
   365 => x"06705651",
   366 => x"5372802e",
   367 => x"a8388480",
   368 => x"808aa604",
   369 => x"83ffe080",
   370 => x"08528480",
   371 => x"80a2bc51",
   372 => x"84808082",
   373 => x"f52d7282",
   374 => x"2efed338",
   375 => x"ff135372",
   376 => x"fee73872",
   377 => x"547383ff",
   378 => x"e0800c02",
   379 => x"90050d04",
   380 => x"02f4050d",
   381 => x"810b83ff",
   382 => x"f1a00cd0",
   383 => x"08708f2a",
   384 => x"70810651",
   385 => x"515372f3",
   386 => x"3872d00c",
   387 => x"84808087",
   388 => x"e62d8480",
   389 => x"80a2d851",
   390 => x"84808085",
   391 => x"d72dd008",
   392 => x"708f2a70",
   393 => x"81065151",
   394 => x"5372f338",
   395 => x"810bd00c",
   396 => x"87538052",
   397 => x"84d480c0",
   398 => x"51848080",
   399 => x"86f12d83",
   400 => x"ffe08008",
   401 => x"812e9738",
   402 => x"72822e09",
   403 => x"81068938",
   404 => x"80538480",
   405 => x"808d9804",
   406 => x"ff135372",
   407 => x"d5388480",
   408 => x"8089ba2d",
   409 => x"83ffe080",
   410 => x"0883fff1",
   411 => x"a00c8152",
   412 => x"87fc80d0",
   413 => x"51848080",
   414 => x"86f12d81",
   415 => x"ff0bd40c",
   416 => x"d008708f",
   417 => x"2a708106",
   418 => x"51515372",
   419 => x"f33872d0",
   420 => x"0c81ff0b",
   421 => x"d40c8153",
   422 => x"7283ffe0",
   423 => x"800c028c",
   424 => x"050d0480",
   425 => x"0b83ffe0",
   426 => x"800c0402",
   427 => x"e0050d79",
   428 => x"7b575780",
   429 => x"5881ff0b",
   430 => x"d40cd008",
   431 => x"708f2a70",
   432 => x"81065151",
   433 => x"5473f338",
   434 => x"82810bd0",
   435 => x"0c81ff0b",
   436 => x"d40c7652",
   437 => x"87fc80d1",
   438 => x"51848080",
   439 => x"86f12d80",
   440 => x"dbc6df55",
   441 => x"83ffe080",
   442 => x"08802e9b",
   443 => x"3883ffe0",
   444 => x"80085376",
   445 => x"52848080",
   446 => x"a2e45184",
   447 => x"808082f5",
   448 => x"2d848080",
   449 => x"8edd0481",
   450 => x"ff0bd40c",
   451 => x"d4087081",
   452 => x"ff065154",
   453 => x"7381fe2e",
   454 => x"098106a5",
   455 => x"3880ff54",
   456 => x"84808086",
   457 => x"a12d83ff",
   458 => x"e0800876",
   459 => x"70840558",
   460 => x"0cff1454",
   461 => x"738025e8",
   462 => x"38815884",
   463 => x"80808ec7",
   464 => x"04ff1555",
   465 => x"74c13881",
   466 => x"ff0bd40c",
   467 => x"d008708f",
   468 => x"2a708106",
   469 => x"51515473",
   470 => x"f33873d0",
   471 => x"0c7783ff",
   472 => x"e0800c02",
   473 => x"a0050d04",
   474 => x"02f4050d",
   475 => x"7470882a",
   476 => x"83fe8006",
   477 => x"7072982a",
   478 => x"0772882b",
   479 => x"87fc8080",
   480 => x"0673982b",
   481 => x"81f00a06",
   482 => x"71730707",
   483 => x"83ffe080",
   484 => x"0c565153",
   485 => x"51028c05",
   486 => x"0d0402f8",
   487 => x"050d028e",
   488 => x"05848080",
   489 => x"80f52d74",
   490 => x"882b0770",
   491 => x"83ffff06",
   492 => x"83ffe080",
   493 => x"0c510288",
   494 => x"050d0402",
   495 => x"f8050d73",
   496 => x"70902b71",
   497 => x"902a0783",
   498 => x"ffe0800c",
   499 => x"52028805",
   500 => x"0d0402ec",
   501 => x"050d800b",
   502 => x"fc800c84",
   503 => x"8080a384",
   504 => x"51848080",
   505 => x"85d72d84",
   506 => x"80808bf0",
   507 => x"2d83ffe0",
   508 => x"8008802e",
   509 => x"82863884",
   510 => x"8080a39c",
   511 => x"51848080",
   512 => x"85d72d84",
   513 => x"808092e0",
   514 => x"2d83ffe1",
   515 => x"a0528480",
   516 => x"80a3b451",
   517 => x"848080a0",
   518 => x"b32d83ff",
   519 => x"e0800880",
   520 => x"2e81cd38",
   521 => x"83ffe1a0",
   522 => x"0b848080",
   523 => x"a3c05254",
   524 => x"84808085",
   525 => x"d72d8055",
   526 => x"73708105",
   527 => x"55848080",
   528 => x"80f52d53",
   529 => x"72a02e80",
   530 => x"e63872c0",
   531 => x"0c72a32e",
   532 => x"81843872",
   533 => x"80c72e09",
   534 => x"81068d38",
   535 => x"84808080",
   536 => x"922d8480",
   537 => x"80918a04",
   538 => x"728a2e09",
   539 => x"81068d38",
   540 => x"84808080",
   541 => x"8c2d8480",
   542 => x"80918a04",
   543 => x"7280cc2e",
   544 => x"09810686",
   545 => x"3883ffe1",
   546 => x"a0547281",
   547 => x"df06f005",
   548 => x"7081ff06",
   549 => x"5153b873",
   550 => x"278938ef",
   551 => x"137081ff",
   552 => x"06515374",
   553 => x"842b7307",
   554 => x"55848080",
   555 => x"90b80472",
   556 => x"a32ea338",
   557 => x"73708105",
   558 => x"55848080",
   559 => x"80f52d53",
   560 => x"72a02ef0",
   561 => x"38ff1475",
   562 => x"53705254",
   563 => x"848080a0",
   564 => x"b32d74fc",
   565 => x"800c7370",
   566 => x"81055584",
   567 => x"808080f5",
   568 => x"2d53728a",
   569 => x"2e098106",
   570 => x"ed388480",
   571 => x"8090b604",
   572 => x"848080a3",
   573 => x"d4518480",
   574 => x"8085d72d",
   575 => x"848080a3",
   576 => x"f0518480",
   577 => x"8085d72d",
   578 => x"800b83ff",
   579 => x"e0800c02",
   580 => x"94050d04",
   581 => x"02e8050d",
   582 => x"77797b58",
   583 => x"55558053",
   584 => x"727625af",
   585 => x"38747081",
   586 => x"05568480",
   587 => x"8080f52d",
   588 => x"74708105",
   589 => x"56848080",
   590 => x"80f52d52",
   591 => x"5271712e",
   592 => x"89388151",
   593 => x"84808092",
   594 => x"d5048113",
   595 => x"53848080",
   596 => x"92a00480",
   597 => x"517083ff",
   598 => x"e0800c02",
   599 => x"98050d04",
   600 => x"02d8050d",
   601 => x"800b83ff",
   602 => x"f5dc0c84",
   603 => x"8080a3fc",
   604 => x"51848080",
   605 => x"85d72d83",
   606 => x"fff1b852",
   607 => x"80518480",
   608 => x"808dab2d",
   609 => x"83ffe080",
   610 => x"085483ff",
   611 => x"e0800895",
   612 => x"38848080",
   613 => x"a48c5184",
   614 => x"808085d7",
   615 => x"2d735584",
   616 => x"80809b8f",
   617 => x"04848080",
   618 => x"a4a05184",
   619 => x"808085d7",
   620 => x"2d805681",
   621 => x"0b83fff1",
   622 => x"ac0c8853",
   623 => x"848080a4",
   624 => x"b85283ff",
   625 => x"f1ee5184",
   626 => x"80809294",
   627 => x"2d83ffe0",
   628 => x"8008762e",
   629 => x"0981068b",
   630 => x"3883ffe0",
   631 => x"800883ff",
   632 => x"f1ac0c88",
   633 => x"53848080",
   634 => x"a4c45283",
   635 => x"fff28a51",
   636 => x"84808092",
   637 => x"942d83ff",
   638 => x"e080088b",
   639 => x"3883ffe0",
   640 => x"800883ff",
   641 => x"f1ac0c83",
   642 => x"fff1ac08",
   643 => x"52848080",
   644 => x"a4d05184",
   645 => x"808082f5",
   646 => x"2d83fff1",
   647 => x"ac08802e",
   648 => x"81cb3883",
   649 => x"fff4fe0b",
   650 => x"84808080",
   651 => x"f52d83ff",
   652 => x"f4ff0b84",
   653 => x"808080f5",
   654 => x"2d71982b",
   655 => x"71902b07",
   656 => x"83fff580",
   657 => x"0b848080",
   658 => x"80f52d70",
   659 => x"882b7207",
   660 => x"83fff581",
   661 => x"0b848080",
   662 => x"80f52d71",
   663 => x"0783fff5",
   664 => x"b60b8480",
   665 => x"8080f52d",
   666 => x"83fff5b7",
   667 => x"0b848080",
   668 => x"80f52d71",
   669 => x"882b0753",
   670 => x"5f54525a",
   671 => x"56575573",
   672 => x"81abaa2e",
   673 => x"09810695",
   674 => x"38755184",
   675 => x"80808ee8",
   676 => x"2d83ffe0",
   677 => x"80085684",
   678 => x"808095b6",
   679 => x"047382d4",
   680 => x"d52e9338",
   681 => x"848080a4",
   682 => x"e4518480",
   683 => x"8085d72d",
   684 => x"84808097",
   685 => x"c2047552",
   686 => x"848080a5",
   687 => x"84518480",
   688 => x"8082f52d",
   689 => x"83fff1b8",
   690 => x"52755184",
   691 => x"80808dab",
   692 => x"2d83ffe0",
   693 => x"80085583",
   694 => x"ffe08008",
   695 => x"802e85af",
   696 => x"38848080",
   697 => x"a59c5184",
   698 => x"808085d7",
   699 => x"2d848080",
   700 => x"a5c45184",
   701 => x"808082f5",
   702 => x"2d885384",
   703 => x"8080a4c4",
   704 => x"5283fff2",
   705 => x"8a518480",
   706 => x"8092942d",
   707 => x"83ffe080",
   708 => x"088e3881",
   709 => x"0b83fff5",
   710 => x"dc0c8480",
   711 => x"8096ce04",
   712 => x"88538480",
   713 => x"80a4b852",
   714 => x"83fff1ee",
   715 => x"51848080",
   716 => x"92942d83",
   717 => x"ffe08008",
   718 => x"802e9338",
   719 => x"848080a5",
   720 => x"dc518480",
   721 => x"8082f52d",
   722 => x"84808097",
   723 => x"c20483ff",
   724 => x"f5b60b84",
   725 => x"808080f5",
   726 => x"2d547380",
   727 => x"d52e0981",
   728 => x"0680df38",
   729 => x"83fff5b7",
   730 => x"0b848080",
   731 => x"80f52d54",
   732 => x"7381aa2e",
   733 => x"09810680",
   734 => x"c938800b",
   735 => x"83fff1b8",
   736 => x"0b848080",
   737 => x"80f52d56",
   738 => x"547481e9",
   739 => x"2e833881",
   740 => x"547481eb",
   741 => x"2e8c3880",
   742 => x"5573752e",
   743 => x"09810683",
   744 => x"ee3883ff",
   745 => x"f1c30b84",
   746 => x"808080f5",
   747 => x"2d597892",
   748 => x"3883fff1",
   749 => x"c40b8480",
   750 => x"8080f52d",
   751 => x"5473822e",
   752 => x"89388055",
   753 => x"8480809b",
   754 => x"8f0483ff",
   755 => x"f1c50b84",
   756 => x"808080f5",
   757 => x"2d7083ff",
   758 => x"f5e40cff",
   759 => x"117083ff",
   760 => x"f5d80c54",
   761 => x"52848080",
   762 => x"a5fc5184",
   763 => x"808082f5",
   764 => x"2d83fff1",
   765 => x"c60b8480",
   766 => x"8080f52d",
   767 => x"83fff1c7",
   768 => x"0b848080",
   769 => x"80f52d56",
   770 => x"76057582",
   771 => x"80290570",
   772 => x"83fff5cc",
   773 => x"0c83fff1",
   774 => x"c80b8480",
   775 => x"8080f52d",
   776 => x"7083fff5",
   777 => x"c80c83ff",
   778 => x"f5dc0859",
   779 => x"57587680",
   780 => x"2e81ec38",
   781 => x"88538480",
   782 => x"80a4c452",
   783 => x"83fff28a",
   784 => x"51848080",
   785 => x"92942d78",
   786 => x"5583ffe0",
   787 => x"800882bf",
   788 => x"3883fff5",
   789 => x"e4087084",
   790 => x"2b83fff5",
   791 => x"b80c7083",
   792 => x"fff5e00c",
   793 => x"83fff1dd",
   794 => x"0b848080",
   795 => x"80f52d83",
   796 => x"fff1dc0b",
   797 => x"84808080",
   798 => x"f52d7182",
   799 => x"80290583",
   800 => x"fff1de0b",
   801 => x"84808080",
   802 => x"f52d7084",
   803 => x"80802912",
   804 => x"83fff1df",
   805 => x"0b848080",
   806 => x"80f52d70",
   807 => x"81800a29",
   808 => x"127083ff",
   809 => x"f1b00c83",
   810 => x"fff5c808",
   811 => x"712983ff",
   812 => x"f5cc0805",
   813 => x"7083fff5",
   814 => x"ec0c83ff",
   815 => x"f1e50b84",
   816 => x"808080f5",
   817 => x"2d83fff1",
   818 => x"e40b8480",
   819 => x"8080f52d",
   820 => x"71828029",
   821 => x"0583fff1",
   822 => x"e60b8480",
   823 => x"8080f52d",
   824 => x"70848080",
   825 => x"291283ff",
   826 => x"f1e70b84",
   827 => x"808080f5",
   828 => x"2d70982b",
   829 => x"81f00a06",
   830 => x"72057083",
   831 => x"fff1b40c",
   832 => x"fe117e29",
   833 => x"770583ff",
   834 => x"f5d40c52",
   835 => x"5752575d",
   836 => x"5751525f",
   837 => x"525c5757",
   838 => x"57848080",
   839 => x"9b8d0483",
   840 => x"fff1ca0b",
   841 => x"84808080",
   842 => x"f52d83ff",
   843 => x"f1c90b84",
   844 => x"808080f5",
   845 => x"2d718280",
   846 => x"29057083",
   847 => x"fff5b80c",
   848 => x"70a02983",
   849 => x"ff057089",
   850 => x"2a7083ff",
   851 => x"f5e00c83",
   852 => x"fff1cf0b",
   853 => x"84808080",
   854 => x"f52d83ff",
   855 => x"f1ce0b84",
   856 => x"808080f5",
   857 => x"2d718280",
   858 => x"29057083",
   859 => x"fff1b00c",
   860 => x"7b71291e",
   861 => x"7083fff5",
   862 => x"d40c7d83",
   863 => x"fff1b40c",
   864 => x"730583ff",
   865 => x"f5ec0c55",
   866 => x"5e515155",
   867 => x"55815574",
   868 => x"83ffe080",
   869 => x"0c02a805",
   870 => x"0d0402ec",
   871 => x"050d7670",
   872 => x"872c7180",
   873 => x"ff065755",
   874 => x"5383fff5",
   875 => x"dc088a38",
   876 => x"72882c73",
   877 => x"81ff0656",
   878 => x"5483fff5",
   879 => x"cc081452",
   880 => x"848080a6",
   881 => x"a0518480",
   882 => x"8082f52d",
   883 => x"83fff1b8",
   884 => x"5283fff5",
   885 => x"cc081451",
   886 => x"8480808d",
   887 => x"ab2d83ff",
   888 => x"e0800853",
   889 => x"83ffe080",
   890 => x"08802e80",
   891 => x"c93883ff",
   892 => x"f5dc0880",
   893 => x"2ea23874",
   894 => x"842983ff",
   895 => x"f1b80570",
   896 => x"08525384",
   897 => x"80808ee8",
   898 => x"2d83ffe0",
   899 => x"8008f00a",
   900 => x"06558480",
   901 => x"809cb404",
   902 => x"741083ff",
   903 => x"f1b80570",
   904 => x"84808080",
   905 => x"e02d5253",
   906 => x"8480808f",
   907 => x"9a2d83ff",
   908 => x"e0800855",
   909 => x"74537283",
   910 => x"ffe0800c",
   911 => x"0294050d",
   912 => x"0402c805",
   913 => x"0d7f615f",
   914 => x"5c800b83",
   915 => x"fff1b408",
   916 => x"83fff5d4",
   917 => x"08585957",
   918 => x"83fff5dc",
   919 => x"08772e8f",
   920 => x"3883fff5",
   921 => x"e408842b",
   922 => x"59848080",
   923 => x"9cf70483",
   924 => x"fff5e008",
   925 => x"842b5980",
   926 => x"5a797927",
   927 => x"81dc3879",
   928 => x"8f06a018",
   929 => x"58547396",
   930 => x"3883fff1",
   931 => x"b8527551",
   932 => x"81165684",
   933 => x"80808dab",
   934 => x"2d83fff1",
   935 => x"b8578077",
   936 => x"84808080",
   937 => x"f52d5654",
   938 => x"74742e83",
   939 => x"38815474",
   940 => x"81e52e81",
   941 => x"9c388170",
   942 => x"7506555d",
   943 => x"73802e81",
   944 => x"90388b17",
   945 => x"84808080",
   946 => x"f52d9806",
   947 => x"5b7a8181",
   948 => x"388b537d",
   949 => x"52765184",
   950 => x"80809294",
   951 => x"2d83ffe0",
   952 => x"800880ed",
   953 => x"389c1708",
   954 => x"51848080",
   955 => x"8ee82d83",
   956 => x"ffe08008",
   957 => x"841d0c9a",
   958 => x"17848080",
   959 => x"80e02d51",
   960 => x"8480808f",
   961 => x"9a2d83ff",
   962 => x"e0800883",
   963 => x"ffe08008",
   964 => x"881e0c83",
   965 => x"ffe08008",
   966 => x"555583ff",
   967 => x"f5dc0880",
   968 => x"2ea03894",
   969 => x"17848080",
   970 => x"80e02d51",
   971 => x"8480808f",
   972 => x"9a2d83ff",
   973 => x"e0800890",
   974 => x"2b83fff0",
   975 => x"0a067016",
   976 => x"51547388",
   977 => x"1d0c7a7c",
   978 => x"0c7c5484",
   979 => x"80809fac",
   980 => x"04811a5a",
   981 => x"8480809c",
   982 => x"f90483ff",
   983 => x"f5dc0880",
   984 => x"2e80c738",
   985 => x"77518480",
   986 => x"809b9a2d",
   987 => x"83ffe080",
   988 => x"0883ffe0",
   989 => x"80085384",
   990 => x"8080a6c0",
   991 => x"52588480",
   992 => x"8082f52d",
   993 => x"7780ffff",
   994 => x"fff80654",
   995 => x"7380ffff",
   996 => x"fff82e96",
   997 => x"38fe1883",
   998 => x"fff5e408",
   999 => x"2983fff5",
  1000 => x"ec080556",
  1001 => x"8480809c",
  1002 => x"f7048054",
  1003 => x"7383ffe0",
  1004 => x"800c02b8",
  1005 => x"050d0402",
  1006 => x"f4050d74",
  1007 => x"70088105",
  1008 => x"710c7008",
  1009 => x"83fff5d8",
  1010 => x"08065353",
  1011 => x"71933888",
  1012 => x"13085184",
  1013 => x"80809b9a",
  1014 => x"2d83ffe0",
  1015 => x"80088814",
  1016 => x"0c810b83",
  1017 => x"ffe0800c",
  1018 => x"028c050d",
  1019 => x"0402f005",
  1020 => x"0d758811",
  1021 => x"08fe0583",
  1022 => x"fff5e408",
  1023 => x"2983fff5",
  1024 => x"ec081172",
  1025 => x"0883fff5",
  1026 => x"d8080605",
  1027 => x"79555354",
  1028 => x"54848080",
  1029 => x"8dab2d83",
  1030 => x"ffe08008",
  1031 => x"5383ffe0",
  1032 => x"8008802e",
  1033 => x"83388153",
  1034 => x"7283ffe0",
  1035 => x"800c0290",
  1036 => x"050d0402",
  1037 => x"ec050d76",
  1038 => x"78715483",
  1039 => x"fff5bc53",
  1040 => x"54558480",
  1041 => x"809cc12d",
  1042 => x"83ffe080",
  1043 => x"085483ff",
  1044 => x"e0800880",
  1045 => x"2e80ce38",
  1046 => x"848080a6",
  1047 => x"d8518480",
  1048 => x"8085d72d",
  1049 => x"83fff5c0",
  1050 => x"0883ff05",
  1051 => x"892a5580",
  1052 => x"54737525",
  1053 => x"80d13872",
  1054 => x"5283fff5",
  1055 => x"bc518480",
  1056 => x"809fed2d",
  1057 => x"83ffe080",
  1058 => x"08802eaf",
  1059 => x"3883fff5",
  1060 => x"bc518480",
  1061 => x"809fb72d",
  1062 => x"84801381",
  1063 => x"15555384",
  1064 => x"8080a0f1",
  1065 => x"04745284",
  1066 => x"8080a6f4",
  1067 => x"51848080",
  1068 => x"82f52d73",
  1069 => x"53848080",
  1070 => x"a1c90483",
  1071 => x"ffe08008",
  1072 => x"53848080",
  1073 => x"a1c90481",
  1074 => x"537283ff",
  1075 => x"e0800c02",
  1076 => x"94050d04",
  1077 => x"00ffffff",
  1078 => x"ff00ffff",
  1079 => x"ffff00ff",
  1080 => x"ffffff00",
  1081 => x"436d645f",
  1082 => x"696e6974",
  1083 => x"0a000000",
  1084 => x"636d645f",
  1085 => x"434d4438",
  1086 => x"20726573",
  1087 => x"706f6e73",
  1088 => x"653a2025",
  1089 => x"640a0000",
  1090 => x"434d4438",
  1091 => x"5f342072",
  1092 => x"6573706f",
  1093 => x"6e73653a",
  1094 => x"2025640a",
  1095 => x"00000000",
  1096 => x"53444843",
  1097 => x"20496e69",
  1098 => x"7469616c",
  1099 => x"697a6174",
  1100 => x"696f6e20",
  1101 => x"6572726f",
  1102 => x"72210a00",
  1103 => x"434d4435",
  1104 => x"38202564",
  1105 => x"0a202000",
  1106 => x"434d4435",
  1107 => x"385f3220",
  1108 => x"25640a20",
  1109 => x"20000000",
  1110 => x"53504920",
  1111 => x"496e6974",
  1112 => x"28290a00",
  1113 => x"52656164",
  1114 => x"20636f6d",
  1115 => x"6d616e64",
  1116 => x"20666169",
  1117 => x"6c656420",
  1118 => x"61742025",
  1119 => x"64202825",
  1120 => x"64290a00",
  1121 => x"496e6974",
  1122 => x"69616c69",
  1123 => x"7a696e67",
  1124 => x"20534420",
  1125 => x"63617264",
  1126 => x"0a000000",
  1127 => x"48756e74",
  1128 => x"696e6720",
  1129 => x"666f7220",
  1130 => x"70617274",
  1131 => x"6974696f",
  1132 => x"6e0a0000",
  1133 => x"4d414e49",
  1134 => x"46455354",
  1135 => x"4d535400",
  1136 => x"50617273",
  1137 => x"696e6720",
  1138 => x"6d616e69",
  1139 => x"66657374",
  1140 => x"0a000000",
  1141 => x"4c6f6164",
  1142 => x"696e6720",
  1143 => x"6d616e69",
  1144 => x"66657374",
  1145 => x"20666169",
  1146 => x"6c65640a",
  1147 => x"00000000",
  1148 => x"52657475",
  1149 => x"726e696e",
  1150 => x"670a0000",
  1151 => x"52656164",
  1152 => x"696e6720",
  1153 => x"4d42520a",
  1154 => x"00000000",
  1155 => x"52656164",
  1156 => x"206f6620",
  1157 => x"4d425220",
  1158 => x"6661696c",
  1159 => x"65640a00",
  1160 => x"4d425220",
  1161 => x"73756363",
  1162 => x"65737366",
  1163 => x"756c6c79",
  1164 => x"20726561",
  1165 => x"640a0000",
  1166 => x"46415431",
  1167 => x"36202020",
  1168 => x"00000000",
  1169 => x"46415433",
  1170 => x"32202020",
  1171 => x"00000000",
  1172 => x"50617274",
  1173 => x"6974696f",
  1174 => x"6e636f75",
  1175 => x"6e742025",
  1176 => x"640a0000",
  1177 => x"4e6f2070",
  1178 => x"61727469",
  1179 => x"74696f6e",
  1180 => x"20736967",
  1181 => x"6e617475",
  1182 => x"72652066",
  1183 => x"6f756e64",
  1184 => x"0a000000",
  1185 => x"52656164",
  1186 => x"696e6720",
  1187 => x"626f6f74",
  1188 => x"20736563",
  1189 => x"746f7220",
  1190 => x"25640a00",
  1191 => x"52656164",
  1192 => x"20626f6f",
  1193 => x"74207365",
  1194 => x"63746f72",
  1195 => x"2066726f",
  1196 => x"6d206669",
  1197 => x"72737420",
  1198 => x"70617274",
  1199 => x"6974696f",
  1200 => x"6e0a0000",
  1201 => x"48756e74",
  1202 => x"696e6720",
  1203 => x"666f7220",
  1204 => x"66696c65",
  1205 => x"73797374",
  1206 => x"656d0a00",
  1207 => x"556e7375",
  1208 => x"70706f72",
  1209 => x"74656420",
  1210 => x"70617274",
  1211 => x"6974696f",
  1212 => x"6e207479",
  1213 => x"7065210d",
  1214 => x"00000000",
  1215 => x"436c7573",
  1216 => x"74657220",
  1217 => x"73697a65",
  1218 => x"3a202564",
  1219 => x"2c20436c",
  1220 => x"75737465",
  1221 => x"72206d61",
  1222 => x"736b2c20",
  1223 => x"25640a00",
  1224 => x"47657443",
  1225 => x"6c757374",
  1226 => x"65722072",
  1227 => x"65616469",
  1228 => x"6e672073",
  1229 => x"6563746f",
  1230 => x"72202564",
  1231 => x"0a000000",
  1232 => x"47657446",
  1233 => x"41544c69",
  1234 => x"6e6b2072",
  1235 => x"65747572",
  1236 => x"6e656420",
  1237 => x"25640a00",
  1238 => x"4f70656e",
  1239 => x"65642066",
  1240 => x"696c652c",
  1241 => x"206c6f61",
  1242 => x"64696e67",
  1243 => x"2e2e2e0a",
  1244 => x"00000000",
  1245 => x"43616e27",
  1246 => x"74206f70",
  1247 => x"656e2025",
  1248 => x"730a0000",
	others => x"00000000"
);

begin

process (clk)
begin
	if (clk'event and clk = '1') then
		if (from_zpu.memAWriteEnable = '1') and (from_zpu.memBWriteEnable = '1') and (from_zpu.memAAddr=from_zpu.memBAddr) and (from_zpu.memAWrite/=from_zpu.memBWrite) then
			report "write collision" severity failure;
		end if;
	
		if (from_zpu.memAWriteEnable = '1') then
			ram(to_integer(unsigned(from_zpu.memAAddr(maxAddrBitBRAM downto 2)))) := from_zpu.memAWrite;
			to_zpu.memARead <= from_zpu.memAWrite;
		else
			to_zpu.memARead <= ram(to_integer(unsigned(from_zpu.memAAddr(maxAddrBitBRAM downto 2))));
		end if;
	end if;
end process;

process (clk)
begin
	if (clk'event and clk = '1') then
		if (from_zpu.memBWriteEnable = '1') then
			ram(to_integer(unsigned(from_zpu.memBAddr(maxAddrBitBRAM downto 2)))) := from_zpu.memBWrite;
			to_zpu.memBRead <= from_zpu.memBWrite;
		else
			to_zpu.memBRead <= ram(to_integer(unsigned(from_zpu.memBAddr(maxAddrBitBRAM downto 2))));
		end if;
	end if;
end process;


end arch;

