-- ZPU
--
-- Copyright 2004-2008 oharboe - �yvind Harboe - oyvind.harboe@zylin.com
-- Modified by Alastair M. Robinson for the ZPUFlex project.
--
-- The FreeBSD license
-- 
-- Redistribution and use in source and binary forms, with or without
-- modification, are permitted provided that the following conditions
-- are met:
-- 
-- 1. Redistributions of source code must retain the above copyright
--    notice, this list of conditions and the following disclaimer.
-- 2. Redistributions in binary form must reproduce the above
--    copyright notice, this list of conditions and the following
--    disclaimer in the documentation and/or other materials
--    provided with the distribution.
-- 
-- THIS SOFTWARE IS PROVIDED BY THE ZPU PROJECT ``AS IS'' AND ANY
-- EXPRESS OR IMPLIED WARRANTIES, INCLUDING, BUT NOT LIMITED TO,
-- THE IMPLIED WARRANTIES OF MERCHANTABILITY AND FITNESS FOR A
-- PARTICULAR PURPOSE ARE DISCLAIMED. IN NO EVENT SHALL THE
-- ZPU PROJECT OR CONTRIBUTORS BE LIABLE FOR ANY DIRECT,
-- INDIRECT, INCIDENTAL, SPECIAL, EXEMPLARY, OR CONSEQUENTIAL DAMAGES
-- (INCLUDING, BUT NOT LIMITED TO, PROCUREMENT OF SUBSTITUTE GOODS
-- OR SERVICES; LOSS OF USE, DATA, OR PROFITS; OR BUSINESS INTERRUPTION)
-- HOWEVER CAUSED AND ON ANY THEORY OF LIABILITY, WHETHER IN CONTRACT,
-- STRICT LIABILITY, OR TORT (INCLUDING NEGLIGENCE OR OTHERWISE)
-- ARISING IN ANY WAY OUT OF THE USE OF THIS SOFTWARE, EVEN IF
-- ADVISED OF THE POSSIBILITY OF SUCH DAMAGE.
-- 
-- The views and conclusions contained in the software and documentation
-- are those of the authors and should not be interpreted as representing
-- official policies, either expressed or implied, of the ZPU Project.

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;


library work;
use work.zpupkg.all;

entity SDBootstrap_ROM is
generic
	(
		maxAddrBitBRAM : integer := maxAddrBitBRAMLimit -- Specify your actual ROM size to save LEs and unnecessary block RAM usage.
	);
port (
	clk : in std_logic;
	areset : in std_logic := '0';
	from_zpu : in ZPU_ToROM;
	to_zpu : out ZPU_FromROM
);
end SDBootstrap_ROM;

architecture arch of SDBootstrap_ROM is

type ram_type is array(natural range 0 to ((2**(maxAddrBitBRAM+1))/4)-1) of std_logic_vector(wordSize-1 downto 0);

shared variable ram : ram_type :=
(
     0 => x"84808080",
     1 => x"8c0b8480",
     2 => x"8081e004",
     3 => x"84808080",
     4 => x"8c04ff0d",
     5 => x"80040400",
     6 => x"40000016",
     7 => x"00000000",
     8 => x"0b83ffe0",
     9 => x"80080b83",
    10 => x"ffe08408",
    11 => x"0b83ffe0",
    12 => x"88088480",
    13 => x"80809808",
    14 => x"2d0b83ff",
    15 => x"e0880c0b",
    16 => x"83ffe084",
    17 => x"0c0b83ff",
    18 => x"e0800c04",
    19 => x"00000000",
    20 => x"00000000",
    21 => x"00000000",
    22 => x"00000000",
    23 => x"00000000",
    24 => x"71fd0608",
    25 => x"72830609",
    26 => x"81058205",
    27 => x"832b2a83",
    28 => x"ffff0652",
    29 => x"0471fc06",
    30 => x"08728306",
    31 => x"09810583",
    32 => x"05101010",
    33 => x"2a81ff06",
    34 => x"520471fd",
    35 => x"060883ff",
    36 => x"ff738306",
    37 => x"09810582",
    38 => x"05832b2b",
    39 => x"09067383",
    40 => x"ffff0673",
    41 => x"83060981",
    42 => x"05820583",
    43 => x"2b0b2b07",
    44 => x"72fc060c",
    45 => x"51510471",
    46 => x"fc060884",
    47 => x"8080a1dc",
    48 => x"73830610",
    49 => x"10050806",
    50 => x"7381ff06",
    51 => x"73830609",
    52 => x"81058305",
    53 => x"1010102b",
    54 => x"0772fc06",
    55 => x"0c515104",
    56 => x"83ffe080",
    57 => x"7083fff5",
    58 => x"f0278e38",
    59 => x"80717084",
    60 => x"05530c84",
    61 => x"808081e4",
    62 => x"04848080",
    63 => x"808c5184",
    64 => x"80808fd9",
    65 => x"0402ec05",
    66 => x"0d765380",
    67 => x"55727525",
    68 => x"8e38ad51",
    69 => x"84808085",
    70 => x"b32d7209",
    71 => x"81055372",
    72 => x"802ebe38",
    73 => x"8754729c",
    74 => x"2a73842b",
    75 => x"54527180",
    76 => x"2e833881",
    77 => x"55897225",
    78 => x"8a38b712",
    79 => x"52848080",
    80 => x"82c604b0",
    81 => x"12527480",
    82 => x"2e893871",
    83 => x"51848080",
    84 => x"85b32dff",
    85 => x"14547380",
    86 => x"25cc3884",
    87 => x"808082e9",
    88 => x"04b05184",
    89 => x"808085b3",
    90 => x"2d800b83",
    91 => x"ffe0800c",
    92 => x"0294050d",
    93 => x"0402c005",
    94 => x"0d0280c4",
    95 => x"05578070",
    96 => x"78708405",
    97 => x"5a087241",
    98 => x"5f5d587c",
    99 => x"7084055e",
   100 => x"085a805b",
   101 => x"79982a7a",
   102 => x"882b5b56",
   103 => x"75893877",
   104 => x"5f848080",
   105 => x"85a7047d",
   106 => x"802e81d3",
   107 => x"38805e75",
   108 => x"80e42e8a",
   109 => x"387580f8",
   110 => x"2e098106",
   111 => x"89387684",
   112 => x"1871085e",
   113 => x"58547580",
   114 => x"e42ea638",
   115 => x"7580e426",
   116 => x"8e387580",
   117 => x"e32e80d9",
   118 => x"38848080",
   119 => x"84bf0475",
   120 => x"80f32eb5",
   121 => x"387580f8",
   122 => x"2e8f3884",
   123 => x"808084bf",
   124 => x"048a5384",
   125 => x"808083fb",
   126 => x"04905383",
   127 => x"ffe0e052",
   128 => x"7b518480",
   129 => x"8082852d",
   130 => x"83ffe080",
   131 => x"0883ffe0",
   132 => x"e05a5584",
   133 => x"808084d8",
   134 => x"04768418",
   135 => x"71087054",
   136 => x"5b585484",
   137 => x"808085d7",
   138 => x"2d805584",
   139 => x"808084d8",
   140 => x"04768418",
   141 => x"71085858",
   142 => x"54848080",
   143 => x"858f04a5",
   144 => x"51848080",
   145 => x"85b32d75",
   146 => x"51848080",
   147 => x"85b32d82",
   148 => x"18588480",
   149 => x"80859a04",
   150 => x"74ff1656",
   151 => x"54807425",
   152 => x"b9387870",
   153 => x"81055a84",
   154 => x"808080f5",
   155 => x"2d705256",
   156 => x"84808085",
   157 => x"b32d8118",
   158 => x"58848080",
   159 => x"84d80475",
   160 => x"a52e0981",
   161 => x"06893881",
   162 => x"5e848080",
   163 => x"859a0475",
   164 => x"51848080",
   165 => x"85b32d81",
   166 => x"1858811b",
   167 => x"5b837b25",
   168 => x"fdf23875",
   169 => x"fde5387e",
   170 => x"83ffe080",
   171 => x"0c0280c0",
   172 => x"050d0402",
   173 => x"f8050d73",
   174 => x"52c00870",
   175 => x"882a7081",
   176 => x"06515151",
   177 => x"70802ef1",
   178 => x"3871c00c",
   179 => x"7183ffe0",
   180 => x"800c0288",
   181 => x"050d0402",
   182 => x"e8050d80",
   183 => x"78575575",
   184 => x"70840557",
   185 => x"08538054",
   186 => x"72982a73",
   187 => x"882b5452",
   188 => x"71802ea2",
   189 => x"38c00870",
   190 => x"882a7081",
   191 => x"06515151",
   192 => x"70802ef1",
   193 => x"3871c00c",
   194 => x"81158115",
   195 => x"55558374",
   196 => x"25d63871",
   197 => x"ca387483",
   198 => x"ffe0800c",
   199 => x"0298050d",
   200 => x"0402f405",
   201 => x"0dd45281",
   202 => x"ff720c71",
   203 => x"085381ff",
   204 => x"720c7288",
   205 => x"2b83fe80",
   206 => x"06720870",
   207 => x"81ff0651",
   208 => x"525381ff",
   209 => x"720c7271",
   210 => x"07882b72",
   211 => x"087081ff",
   212 => x"06515253",
   213 => x"81ff720c",
   214 => x"72710788",
   215 => x"2b720870",
   216 => x"81ff0672",
   217 => x"0783ffe0",
   218 => x"800c5253",
   219 => x"028c050d",
   220 => x"0402f405",
   221 => x"0d747671",
   222 => x"81ff06d4",
   223 => x"0c535383",
   224 => x"fff1a008",
   225 => x"85387189",
   226 => x"2b527198",
   227 => x"2ad40c71",
   228 => x"902a7081",
   229 => x"ff06d40c",
   230 => x"5171882a",
   231 => x"7081ff06",
   232 => x"d40c5171",
   233 => x"81ff06d4",
   234 => x"0c72902a",
   235 => x"7081ff06",
   236 => x"d40c51d4",
   237 => x"087081ff",
   238 => x"06515182",
   239 => x"b8bf5270",
   240 => x"81ff2e09",
   241 => x"81069438",
   242 => x"81ff0bd4",
   243 => x"0cd40870",
   244 => x"81ff06ff",
   245 => x"14545151",
   246 => x"71e53870",
   247 => x"83ffe080",
   248 => x"0c028c05",
   249 => x"0d0402fc",
   250 => x"050d81c7",
   251 => x"5181ff0b",
   252 => x"d40cff11",
   253 => x"51708025",
   254 => x"f4380284",
   255 => x"050d0402",
   256 => x"f0050d84",
   257 => x"808087e6",
   258 => x"2d819c9f",
   259 => x"53805287",
   260 => x"fc80f751",
   261 => x"84808086",
   262 => x"f12d83ff",
   263 => x"e0800854",
   264 => x"83ffe080",
   265 => x"08812e09",
   266 => x"8106ae38",
   267 => x"81ff0bd4",
   268 => x"0c820a52",
   269 => x"849c80e9",
   270 => x"51848080",
   271 => x"86f12d83",
   272 => x"ffe08008",
   273 => x"8e3881ff",
   274 => x"0bd40c73",
   275 => x"53848080",
   276 => x"88e00484",
   277 => x"808087e6",
   278 => x"2dff1353",
   279 => x"72ffae38",
   280 => x"7283ffe0",
   281 => x"800c0290",
   282 => x"050d0402",
   283 => x"f4050d81",
   284 => x"ff0bd40c",
   285 => x"848080a1",
   286 => x"ec518480",
   287 => x"8085d72d",
   288 => x"93538052",
   289 => x"87fc80c1",
   290 => x"51848080",
   291 => x"86f12d83",
   292 => x"ffe08008",
   293 => x"8e3881ff",
   294 => x"0bd40c81",
   295 => x"53848080",
   296 => x"89af0484",
   297 => x"808087e6",
   298 => x"2dff1353",
   299 => x"72d43872",
   300 => x"83ffe080",
   301 => x"0c028c05",
   302 => x"0d0402f0",
   303 => x"050d8480",
   304 => x"8087e62d",
   305 => x"83aa5284",
   306 => x"9c80c851",
   307 => x"84808086",
   308 => x"f12d83ff",
   309 => x"e0800883",
   310 => x"ffe08008",
   311 => x"53848080",
   312 => x"a1f85253",
   313 => x"84808082",
   314 => x"f52d7281",
   315 => x"2e098106",
   316 => x"a9388480",
   317 => x"8086a12d",
   318 => x"83ffe080",
   319 => x"0883ffff",
   320 => x"06537283",
   321 => x"aa2ebb38",
   322 => x"83ffe080",
   323 => x"08528480",
   324 => x"80a29051",
   325 => x"84808082",
   326 => x"f52d8480",
   327 => x"8088eb2d",
   328 => x"8480808a",
   329 => x"ba048154",
   330 => x"8480808b",
   331 => x"e5048480",
   332 => x"80a2a851",
   333 => x"84808082",
   334 => x"f52d8054",
   335 => x"8480808b",
   336 => x"e50481ff",
   337 => x"0bd40cb1",
   338 => x"53848080",
   339 => x"87ff2d83",
   340 => x"ffe08008",
   341 => x"802e80fe",
   342 => x"38805287",
   343 => x"fc80fa51",
   344 => x"84808086",
   345 => x"f12d83ff",
   346 => x"e0800880",
   347 => x"d73883ff",
   348 => x"e0800852",
   349 => x"848080a2",
   350 => x"c4518480",
   351 => x"8082f52d",
   352 => x"81ff0bd4",
   353 => x"0cd40870",
   354 => x"81ff0670",
   355 => x"54848080",
   356 => x"a2d05351",
   357 => x"53848080",
   358 => x"82f52d81",
   359 => x"ff0bd40c",
   360 => x"81ff0bd4",
   361 => x"0c81ff0b",
   362 => x"d40c81ff",
   363 => x"0bd40c72",
   364 => x"862a7081",
   365 => x"06705651",
   366 => x"5372802e",
   367 => x"a8388480",
   368 => x"808aa604",
   369 => x"83ffe080",
   370 => x"08528480",
   371 => x"80a2c451",
   372 => x"84808082",
   373 => x"f52d7282",
   374 => x"2efed338",
   375 => x"ff135372",
   376 => x"fee73872",
   377 => x"547383ff",
   378 => x"e0800c02",
   379 => x"90050d04",
   380 => x"02f4050d",
   381 => x"810b83ff",
   382 => x"f1a00cd0",
   383 => x"08708f2a",
   384 => x"70810651",
   385 => x"515372f3",
   386 => x"3872d00c",
   387 => x"84808087",
   388 => x"e62d8480",
   389 => x"80a2e051",
   390 => x"84808085",
   391 => x"d72dd008",
   392 => x"708f2a70",
   393 => x"81065151",
   394 => x"5372f338",
   395 => x"810bd00c",
   396 => x"87538052",
   397 => x"84d480c0",
   398 => x"51848080",
   399 => x"86f12d83",
   400 => x"ffe08008",
   401 => x"812e9738",
   402 => x"72822e09",
   403 => x"81068938",
   404 => x"80538480",
   405 => x"808d9f04",
   406 => x"ff135372",
   407 => x"d5388480",
   408 => x"8089ba2d",
   409 => x"83ffe080",
   410 => x"0883fff1",
   411 => x"a00c83ff",
   412 => x"e080088e",
   413 => x"38815287",
   414 => x"fc80d051",
   415 => x"84808086",
   416 => x"f12d81ff",
   417 => x"0bd40cd0",
   418 => x"08708f2a",
   419 => x"70810651",
   420 => x"515372f3",
   421 => x"3872d00c",
   422 => x"81ff0bd4",
   423 => x"0c815372",
   424 => x"83ffe080",
   425 => x"0c028c05",
   426 => x"0d04800b",
   427 => x"83ffe080",
   428 => x"0c0402e0",
   429 => x"050d797b",
   430 => x"57578058",
   431 => x"81ff0bd4",
   432 => x"0cd00870",
   433 => x"8f2a7081",
   434 => x"06515154",
   435 => x"73f33882",
   436 => x"810bd00c",
   437 => x"81ff0bd4",
   438 => x"0c765287",
   439 => x"fc80d151",
   440 => x"84808086",
   441 => x"f12d80db",
   442 => x"c6df5583",
   443 => x"ffe08008",
   444 => x"802e9b38",
   445 => x"83ffe080",
   446 => x"08537652",
   447 => x"848080a2",
   448 => x"ec518480",
   449 => x"8082f52d",
   450 => x"8480808e",
   451 => x"e40481ff",
   452 => x"0bd40cd4",
   453 => x"087081ff",
   454 => x"06515473",
   455 => x"81fe2e09",
   456 => x"8106a538",
   457 => x"80ff5484",
   458 => x"808086a1",
   459 => x"2d83ffe0",
   460 => x"80087670",
   461 => x"8405580c",
   462 => x"ff145473",
   463 => x"8025e838",
   464 => x"81588480",
   465 => x"808ece04",
   466 => x"ff155574",
   467 => x"c13881ff",
   468 => x"0bd40cd0",
   469 => x"08708f2a",
   470 => x"70810651",
   471 => x"515473f3",
   472 => x"3873d00c",
   473 => x"7783ffe0",
   474 => x"800c02a0",
   475 => x"050d0402",
   476 => x"f4050d74",
   477 => x"70882a83",
   478 => x"fe800670",
   479 => x"72982a07",
   480 => x"72882b87",
   481 => x"fc808006",
   482 => x"73982b81",
   483 => x"f00a0671",
   484 => x"73070783",
   485 => x"ffe0800c",
   486 => x"56515351",
   487 => x"028c050d",
   488 => x"0402f805",
   489 => x"0d028e05",
   490 => x"84808080",
   491 => x"f52d7488",
   492 => x"2b077083",
   493 => x"ffff0683",
   494 => x"ffe0800c",
   495 => x"51028805",
   496 => x"0d0402f8",
   497 => x"050d7370",
   498 => x"902b7190",
   499 => x"2a0783ff",
   500 => x"e0800c52",
   501 => x"0288050d",
   502 => x"0402ec05",
   503 => x"0d800bfc",
   504 => x"800c8480",
   505 => x"80a38c51",
   506 => x"84808085",
   507 => x"d72d8480",
   508 => x"808bf02d",
   509 => x"83ffe080",
   510 => x"08802e82",
   511 => x"86388480",
   512 => x"80a3a451",
   513 => x"84808085",
   514 => x"d72d8480",
   515 => x"8092e72d",
   516 => x"83ffe1a0",
   517 => x"52848080",
   518 => x"a3bc5184",
   519 => x"8080a0ba",
   520 => x"2d83ffe0",
   521 => x"8008802e",
   522 => x"81cd3883",
   523 => x"ffe1a00b",
   524 => x"848080a3",
   525 => x"c8525484",
   526 => x"808085d7",
   527 => x"2d805573",
   528 => x"70810555",
   529 => x"84808080",
   530 => x"f52d5372",
   531 => x"a02e80e6",
   532 => x"3872c00c",
   533 => x"72a32e81",
   534 => x"84387280",
   535 => x"c72e0981",
   536 => x"068d3884",
   537 => x"80808092",
   538 => x"2d848080",
   539 => x"91910472",
   540 => x"8a2e0981",
   541 => x"068d3884",
   542 => x"8080808c",
   543 => x"2d848080",
   544 => x"91910472",
   545 => x"80cc2e09",
   546 => x"81068638",
   547 => x"83ffe1a0",
   548 => x"547281df",
   549 => x"06f00570",
   550 => x"81ff0651",
   551 => x"53b87327",
   552 => x"8938ef13",
   553 => x"7081ff06",
   554 => x"51537484",
   555 => x"2b730755",
   556 => x"84808090",
   557 => x"bf0472a3",
   558 => x"2ea33873",
   559 => x"70810555",
   560 => x"84808080",
   561 => x"f52d5372",
   562 => x"a02ef038",
   563 => x"ff147553",
   564 => x"70525484",
   565 => x"8080a0ba",
   566 => x"2d74fc80",
   567 => x"0c737081",
   568 => x"05558480",
   569 => x"8080f52d",
   570 => x"53728a2e",
   571 => x"098106ed",
   572 => x"38848080",
   573 => x"90bd0484",
   574 => x"8080a3dc",
   575 => x"51848080",
   576 => x"85d72d84",
   577 => x"8080a3f8",
   578 => x"51848080",
   579 => x"85d72d80",
   580 => x"0b83ffe0",
   581 => x"800c0294",
   582 => x"050d0402",
   583 => x"e8050d77",
   584 => x"797b5855",
   585 => x"55805372",
   586 => x"7625af38",
   587 => x"74708105",
   588 => x"56848080",
   589 => x"80f52d74",
   590 => x"70810556",
   591 => x"84808080",
   592 => x"f52d5252",
   593 => x"71712e89",
   594 => x"38815184",
   595 => x"808092dc",
   596 => x"04811353",
   597 => x"84808092",
   598 => x"a7048051",
   599 => x"7083ffe0",
   600 => x"800c0298",
   601 => x"050d0402",
   602 => x"d8050d80",
   603 => x"0b83fff5",
   604 => x"dc0c8480",
   605 => x"80a48451",
   606 => x"84808085",
   607 => x"d72d83ff",
   608 => x"f1b85280",
   609 => x"51848080",
   610 => x"8db22d83",
   611 => x"ffe08008",
   612 => x"5483ffe0",
   613 => x"80089538",
   614 => x"848080a4",
   615 => x"94518480",
   616 => x"8085d72d",
   617 => x"73558480",
   618 => x"809b9604",
   619 => x"848080a4",
   620 => x"a8518480",
   621 => x"8085d72d",
   622 => x"8056810b",
   623 => x"83fff1ac",
   624 => x"0c885384",
   625 => x"8080a4c0",
   626 => x"5283fff1",
   627 => x"ee518480",
   628 => x"80929b2d",
   629 => x"83ffe080",
   630 => x"08762e09",
   631 => x"81068b38",
   632 => x"83ffe080",
   633 => x"0883fff1",
   634 => x"ac0c8853",
   635 => x"848080a4",
   636 => x"cc5283ff",
   637 => x"f28a5184",
   638 => x"8080929b",
   639 => x"2d83ffe0",
   640 => x"80088b38",
   641 => x"83ffe080",
   642 => x"0883fff1",
   643 => x"ac0c83ff",
   644 => x"f1ac0852",
   645 => x"848080a4",
   646 => x"d8518480",
   647 => x"8082f52d",
   648 => x"83fff1ac",
   649 => x"08802e81",
   650 => x"cb3883ff",
   651 => x"f4fe0b84",
   652 => x"808080f5",
   653 => x"2d83fff4",
   654 => x"ff0b8480",
   655 => x"8080f52d",
   656 => x"71982b71",
   657 => x"902b0783",
   658 => x"fff5800b",
   659 => x"84808080",
   660 => x"f52d7088",
   661 => x"2b720783",
   662 => x"fff5810b",
   663 => x"84808080",
   664 => x"f52d7107",
   665 => x"83fff5b6",
   666 => x"0b848080",
   667 => x"80f52d83",
   668 => x"fff5b70b",
   669 => x"84808080",
   670 => x"f52d7188",
   671 => x"2b07535f",
   672 => x"54525a56",
   673 => x"57557381",
   674 => x"abaa2e09",
   675 => x"81069538",
   676 => x"75518480",
   677 => x"808eef2d",
   678 => x"83ffe080",
   679 => x"08568480",
   680 => x"8095bd04",
   681 => x"7382d4d5",
   682 => x"2e933884",
   683 => x"8080a4ec",
   684 => x"51848080",
   685 => x"85d72d84",
   686 => x"808097c9",
   687 => x"04755284",
   688 => x"8080a58c",
   689 => x"51848080",
   690 => x"82f52d83",
   691 => x"fff1b852",
   692 => x"75518480",
   693 => x"808db22d",
   694 => x"83ffe080",
   695 => x"085583ff",
   696 => x"e0800880",
   697 => x"2e85af38",
   698 => x"848080a5",
   699 => x"a4518480",
   700 => x"8085d72d",
   701 => x"848080a5",
   702 => x"cc518480",
   703 => x"8082f52d",
   704 => x"88538480",
   705 => x"80a4cc52",
   706 => x"83fff28a",
   707 => x"51848080",
   708 => x"929b2d83",
   709 => x"ffe08008",
   710 => x"8e38810b",
   711 => x"83fff5dc",
   712 => x"0c848080",
   713 => x"96d50488",
   714 => x"53848080",
   715 => x"a4c05283",
   716 => x"fff1ee51",
   717 => x"84808092",
   718 => x"9b2d83ff",
   719 => x"e0800880",
   720 => x"2e933884",
   721 => x"8080a5e4",
   722 => x"51848080",
   723 => x"82f52d84",
   724 => x"808097c9",
   725 => x"0483fff5",
   726 => x"b60b8480",
   727 => x"8080f52d",
   728 => x"547380d5",
   729 => x"2e098106",
   730 => x"80df3883",
   731 => x"fff5b70b",
   732 => x"84808080",
   733 => x"f52d5473",
   734 => x"81aa2e09",
   735 => x"810680c9",
   736 => x"38800b83",
   737 => x"fff1b80b",
   738 => x"84808080",
   739 => x"f52d5654",
   740 => x"7481e92e",
   741 => x"83388154",
   742 => x"7481eb2e",
   743 => x"8c388055",
   744 => x"73752e09",
   745 => x"810683ee",
   746 => x"3883fff1",
   747 => x"c30b8480",
   748 => x"8080f52d",
   749 => x"59789238",
   750 => x"83fff1c4",
   751 => x"0b848080",
   752 => x"80f52d54",
   753 => x"73822e89",
   754 => x"38805584",
   755 => x"80809b96",
   756 => x"0483fff1",
   757 => x"c50b8480",
   758 => x"8080f52d",
   759 => x"7083fff5",
   760 => x"e40cff11",
   761 => x"7083fff5",
   762 => x"d80c5452",
   763 => x"848080a6",
   764 => x"84518480",
   765 => x"8082f52d",
   766 => x"83fff1c6",
   767 => x"0b848080",
   768 => x"80f52d83",
   769 => x"fff1c70b",
   770 => x"84808080",
   771 => x"f52d5676",
   772 => x"05758280",
   773 => x"29057083",
   774 => x"fff5cc0c",
   775 => x"83fff1c8",
   776 => x"0b848080",
   777 => x"80f52d70",
   778 => x"83fff5c8",
   779 => x"0c83fff5",
   780 => x"dc085957",
   781 => x"5876802e",
   782 => x"81ec3888",
   783 => x"53848080",
   784 => x"a4cc5283",
   785 => x"fff28a51",
   786 => x"84808092",
   787 => x"9b2d7855",
   788 => x"83ffe080",
   789 => x"0882bf38",
   790 => x"83fff5e4",
   791 => x"0870842b",
   792 => x"83fff5b8",
   793 => x"0c7083ff",
   794 => x"f5e00c83",
   795 => x"fff1dd0b",
   796 => x"84808080",
   797 => x"f52d83ff",
   798 => x"f1dc0b84",
   799 => x"808080f5",
   800 => x"2d718280",
   801 => x"290583ff",
   802 => x"f1de0b84",
   803 => x"808080f5",
   804 => x"2d708480",
   805 => x"80291283",
   806 => x"fff1df0b",
   807 => x"84808080",
   808 => x"f52d7081",
   809 => x"800a2912",
   810 => x"7083fff1",
   811 => x"b00c83ff",
   812 => x"f5c80871",
   813 => x"2983fff5",
   814 => x"cc080570",
   815 => x"83fff5ec",
   816 => x"0c83fff1",
   817 => x"e50b8480",
   818 => x"8080f52d",
   819 => x"83fff1e4",
   820 => x"0b848080",
   821 => x"80f52d71",
   822 => x"82802905",
   823 => x"83fff1e6",
   824 => x"0b848080",
   825 => x"80f52d70",
   826 => x"84808029",
   827 => x"1283fff1",
   828 => x"e70b8480",
   829 => x"8080f52d",
   830 => x"70982b81",
   831 => x"f00a0672",
   832 => x"057083ff",
   833 => x"f1b40cfe",
   834 => x"117e2977",
   835 => x"0583fff5",
   836 => x"d40c5257",
   837 => x"52575d57",
   838 => x"51525f52",
   839 => x"5c575757",
   840 => x"8480809b",
   841 => x"940483ff",
   842 => x"f1ca0b84",
   843 => x"808080f5",
   844 => x"2d83fff1",
   845 => x"c90b8480",
   846 => x"8080f52d",
   847 => x"71828029",
   848 => x"057083ff",
   849 => x"f5b80c70",
   850 => x"a02983ff",
   851 => x"0570892a",
   852 => x"7083fff5",
   853 => x"e00c83ff",
   854 => x"f1cf0b84",
   855 => x"808080f5",
   856 => x"2d83fff1",
   857 => x"ce0b8480",
   858 => x"8080f52d",
   859 => x"71828029",
   860 => x"057083ff",
   861 => x"f1b00c7b",
   862 => x"71291e70",
   863 => x"83fff5d4",
   864 => x"0c7d83ff",
   865 => x"f1b40c73",
   866 => x"0583fff5",
   867 => x"ec0c555e",
   868 => x"51515555",
   869 => x"81557483",
   870 => x"ffe0800c",
   871 => x"02a8050d",
   872 => x"0402ec05",
   873 => x"0d767087",
   874 => x"2c7180ff",
   875 => x"06575553",
   876 => x"83fff5dc",
   877 => x"088a3872",
   878 => x"882c7381",
   879 => x"ff065654",
   880 => x"83fff5cc",
   881 => x"08145284",
   882 => x"8080a6a8",
   883 => x"51848080",
   884 => x"82f52d83",
   885 => x"fff1b852",
   886 => x"83fff5cc",
   887 => x"08145184",
   888 => x"80808db2",
   889 => x"2d83ffe0",
   890 => x"80085383",
   891 => x"ffe08008",
   892 => x"802e80c9",
   893 => x"3883fff5",
   894 => x"dc08802e",
   895 => x"a2387484",
   896 => x"2983fff1",
   897 => x"b8057008",
   898 => x"52538480",
   899 => x"808eef2d",
   900 => x"83ffe080",
   901 => x"08f00a06",
   902 => x"55848080",
   903 => x"9cbb0474",
   904 => x"1083fff1",
   905 => x"b8057084",
   906 => x"808080e0",
   907 => x"2d525384",
   908 => x"80808fa1",
   909 => x"2d83ffe0",
   910 => x"80085574",
   911 => x"537283ff",
   912 => x"e0800c02",
   913 => x"94050d04",
   914 => x"02c8050d",
   915 => x"7f615f5c",
   916 => x"800b83ff",
   917 => x"f1b40883",
   918 => x"fff5d408",
   919 => x"58595783",
   920 => x"fff5dc08",
   921 => x"772e8f38",
   922 => x"83fff5e4",
   923 => x"08842b59",
   924 => x"8480809c",
   925 => x"fe0483ff",
   926 => x"f5e00884",
   927 => x"2b59805a",
   928 => x"79792781",
   929 => x"dc38798f",
   930 => x"06a01858",
   931 => x"54739638",
   932 => x"83fff1b8",
   933 => x"52755181",
   934 => x"16568480",
   935 => x"808db22d",
   936 => x"83fff1b8",
   937 => x"57807784",
   938 => x"808080f5",
   939 => x"2d565474",
   940 => x"742e8338",
   941 => x"81547481",
   942 => x"e52e819c",
   943 => x"38817075",
   944 => x"06555d73",
   945 => x"802e8190",
   946 => x"388b1784",
   947 => x"808080f5",
   948 => x"2d98065b",
   949 => x"7a818138",
   950 => x"8b537d52",
   951 => x"76518480",
   952 => x"80929b2d",
   953 => x"83ffe080",
   954 => x"0880ed38",
   955 => x"9c170851",
   956 => x"8480808e",
   957 => x"ef2d83ff",
   958 => x"e0800884",
   959 => x"1d0c9a17",
   960 => x"84808080",
   961 => x"e02d5184",
   962 => x"80808fa1",
   963 => x"2d83ffe0",
   964 => x"800883ff",
   965 => x"e0800888",
   966 => x"1e0c83ff",
   967 => x"e0800855",
   968 => x"5583fff5",
   969 => x"dc08802e",
   970 => x"a0389417",
   971 => x"84808080",
   972 => x"e02d5184",
   973 => x"80808fa1",
   974 => x"2d83ffe0",
   975 => x"8008902b",
   976 => x"83fff00a",
   977 => x"06701651",
   978 => x"5473881d",
   979 => x"0c7a7c0c",
   980 => x"7c548480",
   981 => x"809fb304",
   982 => x"811a5a84",
   983 => x"80809d80",
   984 => x"0483fff5",
   985 => x"dc08802e",
   986 => x"80c73877",
   987 => x"51848080",
   988 => x"9ba12d83",
   989 => x"ffe08008",
   990 => x"83ffe080",
   991 => x"08538480",
   992 => x"80a6c852",
   993 => x"58848080",
   994 => x"82f52d77",
   995 => x"80ffffff",
   996 => x"f8065473",
   997 => x"80ffffff",
   998 => x"f82e9638",
   999 => x"fe1883ff",
  1000 => x"f5e40829",
  1001 => x"83fff5ec",
  1002 => x"08055684",
  1003 => x"80809cfe",
  1004 => x"04805473",
  1005 => x"83ffe080",
  1006 => x"0c02b805",
  1007 => x"0d0402f4",
  1008 => x"050d7470",
  1009 => x"08810571",
  1010 => x"0c700883",
  1011 => x"fff5d808",
  1012 => x"06535371",
  1013 => x"93388813",
  1014 => x"08518480",
  1015 => x"809ba12d",
  1016 => x"83ffe080",
  1017 => x"0888140c",
  1018 => x"810b83ff",
  1019 => x"e0800c02",
  1020 => x"8c050d04",
  1021 => x"02f0050d",
  1022 => x"75881108",
  1023 => x"fe0583ff",
  1024 => x"f5e40829",
  1025 => x"83fff5ec",
  1026 => x"08117208",
  1027 => x"83fff5d8",
  1028 => x"08060579",
  1029 => x"55535454",
  1030 => x"8480808d",
  1031 => x"b22d83ff",
  1032 => x"e0800853",
  1033 => x"83ffe080",
  1034 => x"08802e83",
  1035 => x"38815372",
  1036 => x"83ffe080",
  1037 => x"0c029005",
  1038 => x"0d0402ec",
  1039 => x"050d7678",
  1040 => x"715483ff",
  1041 => x"f5bc5354",
  1042 => x"55848080",
  1043 => x"9cc82d83",
  1044 => x"ffe08008",
  1045 => x"5483ffe0",
  1046 => x"8008802e",
  1047 => x"80ce3884",
  1048 => x"8080a6e0",
  1049 => x"51848080",
  1050 => x"85d72d83",
  1051 => x"fff5c008",
  1052 => x"83ff0589",
  1053 => x"2a558054",
  1054 => x"73752580",
  1055 => x"d1387252",
  1056 => x"83fff5bc",
  1057 => x"51848080",
  1058 => x"9ff42d83",
  1059 => x"ffe08008",
  1060 => x"802eaf38",
  1061 => x"83fff5bc",
  1062 => x"51848080",
  1063 => x"9fbe2d84",
  1064 => x"80138115",
  1065 => x"55538480",
  1066 => x"80a0f804",
  1067 => x"74528480",
  1068 => x"80a6fc51",
  1069 => x"84808082",
  1070 => x"f52d7353",
  1071 => x"848080a1",
  1072 => x"d00483ff",
  1073 => x"e0800853",
  1074 => x"848080a1",
  1075 => x"d0048153",
  1076 => x"7283ffe0",
  1077 => x"800c0294",
  1078 => x"050d0400",
  1079 => x"00ffffff",
  1080 => x"ff00ffff",
  1081 => x"ffff00ff",
  1082 => x"ffffff00",
  1083 => x"436d645f",
  1084 => x"696e6974",
  1085 => x"0a000000",
  1086 => x"636d645f",
  1087 => x"434d4438",
  1088 => x"20726573",
  1089 => x"706f6e73",
  1090 => x"653a2025",
  1091 => x"640a0000",
  1092 => x"434d4438",
  1093 => x"5f342072",
  1094 => x"6573706f",
  1095 => x"6e73653a",
  1096 => x"2025640a",
  1097 => x"00000000",
  1098 => x"53444843",
  1099 => x"20496e69",
  1100 => x"7469616c",
  1101 => x"697a6174",
  1102 => x"696f6e20",
  1103 => x"6572726f",
  1104 => x"72210a00",
  1105 => x"434d4435",
  1106 => x"38202564",
  1107 => x"0a202000",
  1108 => x"434d4435",
  1109 => x"385f3220",
  1110 => x"25640a20",
  1111 => x"20000000",
  1112 => x"53504920",
  1113 => x"496e6974",
  1114 => x"28290a00",
  1115 => x"52656164",
  1116 => x"20636f6d",
  1117 => x"6d616e64",
  1118 => x"20666169",
  1119 => x"6c656420",
  1120 => x"61742025",
  1121 => x"64202825",
  1122 => x"64290a00",
  1123 => x"496e6974",
  1124 => x"69616c69",
  1125 => x"7a696e67",
  1126 => x"20534420",
  1127 => x"63617264",
  1128 => x"0a000000",
  1129 => x"48756e74",
  1130 => x"696e6720",
  1131 => x"666f7220",
  1132 => x"70617274",
  1133 => x"6974696f",
  1134 => x"6e0a0000",
  1135 => x"4d414e49",
  1136 => x"46455354",
  1137 => x"4d535400",
  1138 => x"50617273",
  1139 => x"696e6720",
  1140 => x"6d616e69",
  1141 => x"66657374",
  1142 => x"0a000000",
  1143 => x"4c6f6164",
  1144 => x"696e6720",
  1145 => x"6d616e69",
  1146 => x"66657374",
  1147 => x"20666169",
  1148 => x"6c65640a",
  1149 => x"00000000",
  1150 => x"52657475",
  1151 => x"726e696e",
  1152 => x"670a0000",
  1153 => x"52656164",
  1154 => x"696e6720",
  1155 => x"4d42520a",
  1156 => x"00000000",
  1157 => x"52656164",
  1158 => x"206f6620",
  1159 => x"4d425220",
  1160 => x"6661696c",
  1161 => x"65640a00",
  1162 => x"4d425220",
  1163 => x"73756363",
  1164 => x"65737366",
  1165 => x"756c6c79",
  1166 => x"20726561",
  1167 => x"640a0000",
  1168 => x"46415431",
  1169 => x"36202020",
  1170 => x"00000000",
  1171 => x"46415433",
  1172 => x"32202020",
  1173 => x"00000000",
  1174 => x"50617274",
  1175 => x"6974696f",
  1176 => x"6e636f75",
  1177 => x"6e742025",
  1178 => x"640a0000",
  1179 => x"4e6f2070",
  1180 => x"61727469",
  1181 => x"74696f6e",
  1182 => x"20736967",
  1183 => x"6e617475",
  1184 => x"72652066",
  1185 => x"6f756e64",
  1186 => x"0a000000",
  1187 => x"52656164",
  1188 => x"696e6720",
  1189 => x"626f6f74",
  1190 => x"20736563",
  1191 => x"746f7220",
  1192 => x"25640a00",
  1193 => x"52656164",
  1194 => x"20626f6f",
  1195 => x"74207365",
  1196 => x"63746f72",
  1197 => x"2066726f",
  1198 => x"6d206669",
  1199 => x"72737420",
  1200 => x"70617274",
  1201 => x"6974696f",
  1202 => x"6e0a0000",
  1203 => x"48756e74",
  1204 => x"696e6720",
  1205 => x"666f7220",
  1206 => x"66696c65",
  1207 => x"73797374",
  1208 => x"656d0a00",
  1209 => x"556e7375",
  1210 => x"70706f72",
  1211 => x"74656420",
  1212 => x"70617274",
  1213 => x"6974696f",
  1214 => x"6e207479",
  1215 => x"7065210d",
  1216 => x"00000000",
  1217 => x"436c7573",
  1218 => x"74657220",
  1219 => x"73697a65",
  1220 => x"3a202564",
  1221 => x"2c20436c",
  1222 => x"75737465",
  1223 => x"72206d61",
  1224 => x"736b2c20",
  1225 => x"25640a00",
  1226 => x"47657443",
  1227 => x"6c757374",
  1228 => x"65722072",
  1229 => x"65616469",
  1230 => x"6e672073",
  1231 => x"6563746f",
  1232 => x"72202564",
  1233 => x"0a000000",
  1234 => x"47657446",
  1235 => x"41544c69",
  1236 => x"6e6b2072",
  1237 => x"65747572",
  1238 => x"6e656420",
  1239 => x"25640a00",
  1240 => x"4f70656e",
  1241 => x"65642066",
  1242 => x"696c652c",
  1243 => x"206c6f61",
  1244 => x"64696e67",
  1245 => x"2e2e2e0a",
  1246 => x"00000000",
  1247 => x"43616e27",
  1248 => x"74206f70",
  1249 => x"656e2025",
  1250 => x"730a0000",
	others => x"00000000"
);

begin

process (clk)
begin
	if (clk'event and clk = '1') then
		if (from_zpu.memAWriteEnable = '1') and (from_zpu.memBWriteEnable = '1') and (from_zpu.memAAddr=from_zpu.memBAddr) and (from_zpu.memAWrite/=from_zpu.memBWrite) then
			report "write collision" severity failure;
		end if;
	
		if (from_zpu.memAWriteEnable = '1') then
			ram(to_integer(unsigned(from_zpu.memAAddr(maxAddrBitBRAM downto 2)))) := from_zpu.memAWrite;
			to_zpu.memARead <= from_zpu.memAWrite;
		else
			to_zpu.memARead <= ram(to_integer(unsigned(from_zpu.memAAddr(maxAddrBitBRAM downto 2))));
		end if;
	end if;
end process;

process (clk)
begin
	if (clk'event and clk = '1') then
		if (from_zpu.memBWriteEnable = '1') then
			ram(to_integer(unsigned(from_zpu.memBAddr(maxAddrBitBRAM downto 2)))) := from_zpu.memBWrite;
			to_zpu.memBRead <= from_zpu.memBWrite;
		else
			to_zpu.memBRead <= ram(to_integer(unsigned(from_zpu.memBAddr(maxAddrBitBRAM downto 2))));
		end if;
	end if;
end process;


end arch;

