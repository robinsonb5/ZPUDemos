-- ZPU
--
-- Copyright 2004-2008 oharboe - �yvind Harboe - oyvind.harboe@zylin.com
-- Modified by Alastair M. Robinson for the ZPUFlex project.
--
-- The FreeBSD license
-- 
-- Redistribution and use in source and binary forms, with or without
-- modification, are permitted provided that the following conditions
-- are met:
-- 
-- 1. Redistributions of source code must retain the above copyright
--    notice, this list of conditions and the following disclaimer.
-- 2. Redistributions in binary form must reproduce the above
--    copyright notice, this list of conditions and the following
--    disclaimer in the documentation and/or other materials
--    provided with the distribution.
-- 
-- THIS SOFTWARE IS PROVIDED BY THE ZPU PROJECT ``AS IS'' AND ANY
-- EXPRESS OR IMPLIED WARRANTIES, INCLUDING, BUT NOT LIMITED TO,
-- THE IMPLIED WARRANTIES OF MERCHANTABILITY AND FITNESS FOR A
-- PARTICULAR PURPOSE ARE DISCLAIMED. IN NO EVENT SHALL THE
-- ZPU PROJECT OR CONTRIBUTORS BE LIABLE FOR ANY DIRECT,
-- INDIRECT, INCIDENTAL, SPECIAL, EXEMPLARY, OR CONSEQUENTIAL DAMAGES
-- (INCLUDING, BUT NOT LIMITED TO, PROCUREMENT OF SUBSTITUTE GOODS
-- OR SERVICES; LOSS OF USE, DATA, OR PROFITS; OR BUSINESS INTERRUPTION)
-- HOWEVER CAUSED AND ON ANY THEORY OF LIABILITY, WHETHER IN CONTRACT,
-- STRICT LIABILITY, OR TORT (INCLUDING NEGLIGENCE OR OTHERWISE)
-- ARISING IN ANY WAY OUT OF THE USE OF THIS SOFTWARE, EVEN IF
-- ADVISED OF THE POSSIBILITY OF SUCH DAMAGE.
-- 
-- The views and conclusions contained in the software and documentation
-- are those of the authors and should not be interpreted as representing
-- official policies, either expressed or implied, of the ZPU Project.

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;


library work;
use work.zpu_config.all;
use work.zpupkg.all;

entity Dhrystone_fast_ROM is
generic
	(
		maxAddrBit : integer := maxAddrBitBRAMLimit -- Specify your actual ROM size to save LEs and unnecessary block RAM usage.
	);
port (
	clk : in std_logic;
	areset : in std_logic := '0';
	from_zpu : in ZPU_ToROM;
	to_zpu : out ZPU_FromROM
);
end Dhrystone_fast_ROM;

architecture arch of Dhrystone_fast_ROM is

type ram_type is array(natural range 0 to ((2**(maxAddrBit+1))/4)-1) of std_logic_vector(wordSize-1 downto 0);

shared variable ram : ram_type :=
(
     0 => x"0b0b0b88",
     1 => x"dd040000",
     2 => x"00000000",
     3 => x"00000000",
     4 => x"00000000",
     5 => x"00000000",
     6 => x"00000000",
     7 => x"00000000",
     8 => x"88088c08",
     9 => x"90080b0b",
    10 => x"0b88e708",
    11 => x"2d900c8c",
    12 => x"0c880c04",
    13 => x"00000000",
    14 => x"00000000",
    15 => x"00000000",
    16 => x"71fd0608",
    17 => x"72830609",
    18 => x"81058205",
    19 => x"832b2a83",
    20 => x"ffff0652",
    21 => x"04000000",
    22 => x"00000000",
    23 => x"00000000",
    24 => x"71fd0608",
    25 => x"83ffff73",
    26 => x"83060981",
    27 => x"05820583",
    28 => x"2b2b0906",
    29 => x"7383ffff",
    30 => x"0b0b0b0b",
    31 => x"83a50400",
    32 => x"72098105",
    33 => x"72057373",
    34 => x"09060906",
    35 => x"73097306",
    36 => x"070a8106",
    37 => x"53510400",
    38 => x"00000000",
    39 => x"00000000",
    40 => x"72722473",
    41 => x"732e0753",
    42 => x"51040000",
    43 => x"00000000",
    44 => x"00000000",
    45 => x"00000000",
    46 => x"00000000",
    47 => x"00000000",
    48 => x"71737109",
    49 => x"71068106",
    50 => x"09810572",
    51 => x"0a100a72",
    52 => x"0a100a31",
    53 => x"050a8106",
    54 => x"51515351",
    55 => x"04000000",
    56 => x"72722673",
    57 => x"732e0753",
    58 => x"51040000",
    59 => x"00000000",
    60 => x"00000000",
    61 => x"00000000",
    62 => x"00000000",
    63 => x"00000000",
    64 => x"00000000",
    65 => x"00000000",
    66 => x"00000000",
    67 => x"00000000",
    68 => x"00000000",
    69 => x"00000000",
    70 => x"00000000",
    71 => x"00000000",
    72 => x"0b0b0b88",
    73 => x"ba040000",
    74 => x"00000000",
    75 => x"00000000",
    76 => x"00000000",
    77 => x"00000000",
    78 => x"00000000",
    79 => x"00000000",
    80 => x"720a722b",
    81 => x"0a535104",
    82 => x"00000000",
    83 => x"00000000",
    84 => x"00000000",
    85 => x"00000000",
    86 => x"00000000",
    87 => x"00000000",
    88 => x"72729f06",
    89 => x"0981050b",
    90 => x"0b0b889f",
    91 => x"05040000",
    92 => x"00000000",
    93 => x"00000000",
    94 => x"00000000",
    95 => x"00000000",
    96 => x"72722aff",
    97 => x"739f062a",
    98 => x"0974090a",
    99 => x"8106ff05",
   100 => x"06075351",
   101 => x"04000000",
   102 => x"00000000",
   103 => x"00000000",
   104 => x"71715351",
   105 => x"04067383",
   106 => x"06098105",
   107 => x"8205832b",
   108 => x"0b2b0772",
   109 => x"fc060c51",
   110 => x"51040000",
   111 => x"00000000",
   112 => x"72098105",
   113 => x"72050970",
   114 => x"81050906",
   115 => x"0a810653",
   116 => x"51040000",
   117 => x"00000000",
   118 => x"00000000",
   119 => x"00000000",
   120 => x"72098105",
   121 => x"72050970",
   122 => x"81050906",
   123 => x"0a098106",
   124 => x"53510400",
   125 => x"00000000",
   126 => x"00000000",
   127 => x"00000000",
   128 => x"71098105",
   129 => x"52040000",
   130 => x"00000000",
   131 => x"00000000",
   132 => x"00000000",
   133 => x"00000000",
   134 => x"00000000",
   135 => x"00000000",
   136 => x"72720981",
   137 => x"05055351",
   138 => x"04000000",
   139 => x"00000000",
   140 => x"00000000",
   141 => x"00000000",
   142 => x"00000000",
   143 => x"00000000",
   144 => x"72097206",
   145 => x"73730906",
   146 => x"07535104",
   147 => x"00000000",
   148 => x"00000000",
   149 => x"00000000",
   150 => x"00000000",
   151 => x"00000000",
   152 => x"71fc0608",
   153 => x"72830609",
   154 => x"81058305",
   155 => x"1010102a",
   156 => x"81ff0652",
   157 => x"04000000",
   158 => x"00000000",
   159 => x"00000000",
   160 => x"71fc0608",
   161 => x"0b0b0ba1",
   162 => x"94738306",
   163 => x"10100508",
   164 => x"060b0b0b",
   165 => x"88a20400",
   166 => x"00000000",
   167 => x"00000000",
   168 => x"88088c08",
   169 => x"90087575",
   170 => x"0b0b0b9a",
   171 => x"872d5050",
   172 => x"88085690",
   173 => x"0c8c0c88",
   174 => x"0c510400",
   175 => x"00000000",
   176 => x"88088c08",
   177 => x"90087575",
   178 => x"0b0b0b9b",
   179 => x"b92d5050",
   180 => x"88085690",
   181 => x"0c8c0c88",
   182 => x"0c510400",
   183 => x"00000000",
   184 => x"72097081",
   185 => x"0509060a",
   186 => x"8106ff05",
   187 => x"70547106",
   188 => x"73097274",
   189 => x"05ff0506",
   190 => x"07515151",
   191 => x"04000000",
   192 => x"72097081",
   193 => x"0509060a",
   194 => x"098106ff",
   195 => x"05705471",
   196 => x"06730972",
   197 => x"7405ff05",
   198 => x"06075151",
   199 => x"51040000",
   200 => x"05ff0504",
   201 => x"00000000",
   202 => x"00000000",
   203 => x"00000000",
   204 => x"00000000",
   205 => x"00000000",
   206 => x"00000000",
   207 => x"00000000",
   208 => x"04000000",
   209 => x"00000000",
   210 => x"00000000",
   211 => x"00000000",
   212 => x"00000000",
   213 => x"00000000",
   214 => x"00000000",
   215 => x"00000000",
   216 => x"71810552",
   217 => x"04000000",
   218 => x"00000000",
   219 => x"00000000",
   220 => x"00000000",
   221 => x"00000000",
   222 => x"00000000",
   223 => x"00000000",
   224 => x"00000000",
   225 => x"00000000",
   226 => x"00000000",
   227 => x"00000000",
   228 => x"00000000",
   229 => x"00000000",
   230 => x"00000000",
   231 => x"00000000",
   232 => x"02840572",
   233 => x"10100552",
   234 => x"04000000",
   235 => x"00000000",
   236 => x"00000000",
   237 => x"00000000",
   238 => x"00000000",
   239 => x"00000000",
   240 => x"00000000",
   241 => x"00000000",
   242 => x"00000000",
   243 => x"00000000",
   244 => x"00000000",
   245 => x"00000000",
   246 => x"00000000",
   247 => x"00000000",
   248 => x"717105ff",
   249 => x"05715351",
   250 => x"020d0400",
   251 => x"00000000",
   252 => x"00000000",
   253 => x"00000000",
   254 => x"00000000",
   255 => x"00000000",
   256 => x"10101010",
   257 => x"10101010",
   258 => x"10101010",
   259 => x"10101010",
   260 => x"10101010",
   261 => x"10101010",
   262 => x"10101010",
   263 => x"10101053",
   264 => x"51047381",
   265 => x"ff067383",
   266 => x"06098105",
   267 => x"83051010",
   268 => x"102b0772",
   269 => x"fc060c51",
   270 => x"51047272",
   271 => x"80728106",
   272 => x"ff050972",
   273 => x"06057110",
   274 => x"52720a10",
   275 => x"0a5372ed",
   276 => x"38515153",
   277 => x"51040000",
   278 => x"800488da",
   279 => x"0488da0b",
   280 => x"8fb50404",
   281 => x"00000000",
   282 => x"00046302",
   283 => x"c0050d02",
   284 => x"80c4050b",
   285 => x"0b0ba6bc",
   286 => x"5a5c807c",
   287 => x"7084055e",
   288 => x"08715f5f",
   289 => x"577d7084",
   290 => x"055f0856",
   291 => x"80587598",
   292 => x"2a76882b",
   293 => x"57557480",
   294 => x"2e82d038",
   295 => x"7c802eb9",
   296 => x"38805d74",
   297 => x"80e42e81",
   298 => x"9f387480",
   299 => x"e42680dc",
   300 => x"387480e3",
   301 => x"2eba38a5",
   302 => x"518bf42d",
   303 => x"74518bf4",
   304 => x"2d821757",
   305 => x"81185883",
   306 => x"7825c338",
   307 => x"74ffb638",
   308 => x"7e880c02",
   309 => x"80c0050d",
   310 => x"0474a52e",
   311 => x"09810698",
   312 => x"38810b81",
   313 => x"19595d83",
   314 => x"7825ffa2",
   315 => x"3889cc04",
   316 => x"7b841d71",
   317 => x"08575d5a",
   318 => x"74518bf4",
   319 => x"2d811781",
   320 => x"19595783",
   321 => x"7825ff86",
   322 => x"3889cc04",
   323 => x"7480f32e",
   324 => x"098106ff",
   325 => x"a2387b84",
   326 => x"1d710870",
   327 => x"545b5d54",
   328 => x"8c952d80",
   329 => x"0bff1155",
   330 => x"53807325",
   331 => x"ff963878",
   332 => x"7081055a",
   333 => x"84e02d70",
   334 => x"52558bf4",
   335 => x"2d811774",
   336 => x"ff165654",
   337 => x"578aa904",
   338 => x"7b841d71",
   339 => x"080b0b0b",
   340 => x"a6bc0b0b",
   341 => x"0b0ba5ec",
   342 => x"615f585e",
   343 => x"525d5372",
   344 => x"ba38b00b",
   345 => x"0b0b0ba5",
   346 => x"ec0b8580",
   347 => x"2d811454",
   348 => x"ff145473",
   349 => x"84e02d7b",
   350 => x"7081055d",
   351 => x"85802d81",
   352 => x"1a5a730b",
   353 => x"0b0ba5ec",
   354 => x"2e098106",
   355 => x"e338807b",
   356 => x"85802d79",
   357 => x"ff115553",
   358 => x"8aa9048a",
   359 => x"52725199",
   360 => x"e22d8808",
   361 => x"0b0b0ba1",
   362 => x"a40584e0",
   363 => x"2d747081",
   364 => x"05568580",
   365 => x"2d8a5272",
   366 => x"5199bd2d",
   367 => x"88085388",
   368 => x"08d93873",
   369 => x"0b0b0ba5",
   370 => x"ec2ec338",
   371 => x"ff145473",
   372 => x"84e02d7b",
   373 => x"7081055d",
   374 => x"85802d81",
   375 => x"1a5a730b",
   376 => x"0b0ba5ec",
   377 => x"2effa738",
   378 => x"8af00476",
   379 => x"880c0280",
   380 => x"c0050d04",
   381 => x"02f8050d",
   382 => x"7352c008",
   383 => x"70882a70",
   384 => x"81065151",
   385 => x"5170802e",
   386 => x"f13871c0",
   387 => x"0c71880c",
   388 => x"0288050d",
   389 => x"0402e805",
   390 => x"0d775675",
   391 => x"70840557",
   392 => x"08538054",
   393 => x"72982a73",
   394 => x"882b5452",
   395 => x"71802ea2",
   396 => x"38c00870",
   397 => x"882a7081",
   398 => x"06515151",
   399 => x"70802ef1",
   400 => x"3871c00c",
   401 => x"81158115",
   402 => x"55558374",
   403 => x"25d63871",
   404 => x"ca387488",
   405 => x"0c029805",
   406 => x"0d04c808",
   407 => x"880c0402",
   408 => x"fc050d80",
   409 => x"c10b80f6",
   410 => x"880b8580",
   411 => x"2d800b80",
   412 => x"f8a00c70",
   413 => x"880c0284",
   414 => x"050d0402",
   415 => x"f8050d80",
   416 => x"0b80f688",
   417 => x"0b84e02d",
   418 => x"52527080",
   419 => x"c12e9d38",
   420 => x"7180f8a0",
   421 => x"080780f8",
   422 => x"a00c80c2",
   423 => x"0b80f68c",
   424 => x"0b85802d",
   425 => x"70880c02",
   426 => x"88050d04",
   427 => x"810b80f8",
   428 => x"a0080780",
   429 => x"f8a00c80",
   430 => x"c20b80f6",
   431 => x"8c0b8580",
   432 => x"2d70880c",
   433 => x"0288050d",
   434 => x"0402f005",
   435 => x"0d757008",
   436 => x"8a055353",
   437 => x"80f6880b",
   438 => x"84e02d51",
   439 => x"7080c12e",
   440 => x"8c3873f0",
   441 => x"3870880c",
   442 => x"0290050d",
   443 => x"04ff1270",
   444 => x"80f68408",
   445 => x"31740c88",
   446 => x"0c029005",
   447 => x"0d0402ec",
   448 => x"050d80f6",
   449 => x"b0085574",
   450 => x"802e8c38",
   451 => x"76750871",
   452 => x"0c80f6b0",
   453 => x"0856548c",
   454 => x"155380f6",
   455 => x"8408528a",
   456 => x"5197932d",
   457 => x"73880c02",
   458 => x"94050d04",
   459 => x"02e8050d",
   460 => x"77700856",
   461 => x"56b05380",
   462 => x"f6b00852",
   463 => x"74519ee5",
   464 => x"2d850b8c",
   465 => x"170c850b",
   466 => x"8c160c75",
   467 => x"08750c80",
   468 => x"f6b00854",
   469 => x"73802e8a",
   470 => x"38730875",
   471 => x"0c80f6b0",
   472 => x"08548c14",
   473 => x"5380f684",
   474 => x"08528a51",
   475 => x"97932d84",
   476 => x"1508ae38",
   477 => x"860b8c16",
   478 => x"0c881552",
   479 => x"88160851",
   480 => x"96ad2d80",
   481 => x"f6b00870",
   482 => x"08760c54",
   483 => x"8c157054",
   484 => x"548a5273",
   485 => x"08519793",
   486 => x"2d73880c",
   487 => x"0298050d",
   488 => x"04750854",
   489 => x"b0537352",
   490 => x"75519ee5",
   491 => x"2d73880c",
   492 => x"0298050d",
   493 => x"0402c805",
   494 => x"0d80f59c",
   495 => x"0b80f5d0",
   496 => x"0c80f5d4",
   497 => x"0b80f6b0",
   498 => x"0c80f59c",
   499 => x"0b80f5d4",
   500 => x"0c800b80",
   501 => x"f5d40b84",
   502 => x"050c820b",
   503 => x"80f5d40b",
   504 => x"88050ca8",
   505 => x"0b80f5d4",
   506 => x"0b8c050c",
   507 => x"9f53a1b8",
   508 => x"5280f5e4",
   509 => x"519ee52d",
   510 => x"9f53a1d8",
   511 => x"5280f880",
   512 => x"519ee52d",
   513 => x"8a0bb3e8",
   514 => x"0ca4b851",
   515 => x"88eb2da1",
   516 => x"f85188eb",
   517 => x"2da4b851",
   518 => x"88eb2da5",
   519 => x"e808802e",
   520 => x"849138a2",
   521 => x"a85188eb",
   522 => x"2da4b851",
   523 => x"88eb2da5",
   524 => x"e40852a2",
   525 => x"d45188eb",
   526 => x"2dc80870",
   527 => x"a7880c56",
   528 => x"8158800b",
   529 => x"a5e40825",
   530 => x"82dc3802",
   531 => x"ac055b80",
   532 => x"c10b80f6",
   533 => x"880b8580",
   534 => x"2d810b80",
   535 => x"f8a00c80",
   536 => x"c20b80f6",
   537 => x"8c0b8580",
   538 => x"2d825c83",
   539 => x"5a9f53a3",
   540 => x"845280f6",
   541 => x"90519ee5",
   542 => x"2d815d80",
   543 => x"0b80f690",
   544 => x"5380f880",
   545 => x"525598c5",
   546 => x"2d880875",
   547 => x"2e098106",
   548 => x"83388155",
   549 => x"7480f8a0",
   550 => x"0c7b7057",
   551 => x"55748325",
   552 => x"a1387410",
   553 => x"1015fd05",
   554 => x"5e02b805",
   555 => x"fc055383",
   556 => x"52755197",
   557 => x"932d811c",
   558 => x"705d7057",
   559 => x"55837524",
   560 => x"e1387d54",
   561 => x"7453a78c",
   562 => x"5280f6b8",
   563 => x"5197a52d",
   564 => x"80f6b008",
   565 => x"70085757",
   566 => x"b0537652",
   567 => x"75519ee5",
   568 => x"2d850b8c",
   569 => x"180c850b",
   570 => x"8c170c76",
   571 => x"08760c80",
   572 => x"f6b00855",
   573 => x"74802e8a",
   574 => x"38740876",
   575 => x"0c80f6b0",
   576 => x"08558c15",
   577 => x"5380f684",
   578 => x"08528a51",
   579 => x"97932d84",
   580 => x"160883d8",
   581 => x"38860b8c",
   582 => x"170c8816",
   583 => x"52881708",
   584 => x"5196ad2d",
   585 => x"80f6b008",
   586 => x"7008770c",
   587 => x"578c1670",
   588 => x"54558a52",
   589 => x"74085197",
   590 => x"932d80c1",
   591 => x"0b80f68c",
   592 => x"0b84e02d",
   593 => x"56567575",
   594 => x"26a53880",
   595 => x"c3527551",
   596 => x"98912d88",
   597 => x"087d2e82",
   598 => x"e2388116",
   599 => x"7081ff06",
   600 => x"80f68c0b",
   601 => x"84e02d52",
   602 => x"57557476",
   603 => x"27dd3879",
   604 => x"7c297e53",
   605 => x"519a872d",
   606 => x"88085c88",
   607 => x"088a0580",
   608 => x"f6880b84",
   609 => x"e02d80f6",
   610 => x"84085957",
   611 => x"557580c1",
   612 => x"2e82f438",
   613 => x"78f73881",
   614 => x"1858a5e4",
   615 => x"087825fd",
   616 => x"ae38a788",
   617 => x"0856c808",
   618 => x"7080f5cc",
   619 => x"0c707731",
   620 => x"70a7840c",
   621 => x"53a3a452",
   622 => x"5b88eb2d",
   623 => x"a7840856",
   624 => x"80f77625",
   625 => x"80f338a5",
   626 => x"e4087053",
   627 => x"7687e829",
   628 => x"525a9a87",
   629 => x"2d8808a6",
   630 => x"fc0c7552",
   631 => x"7987e829",
   632 => x"519a872d",
   633 => x"8808a780",
   634 => x"0c755279",
   635 => x"84b92951",
   636 => x"9a872d88",
   637 => x"0880f6b4",
   638 => x"0ca3b451",
   639 => x"88eb2da6",
   640 => x"fc0852a3",
   641 => x"e45188eb",
   642 => x"2da3ec51",
   643 => x"88eb2da7",
   644 => x"800852a3",
   645 => x"e45188eb",
   646 => x"2d80f6b4",
   647 => x"0852a49c",
   648 => x"5188eb2d",
   649 => x"a4b85188",
   650 => x"eb2d800b",
   651 => x"880c02b8",
   652 => x"050d04a4",
   653 => x"bc5190a6",
   654 => x"04a4ec51",
   655 => x"88eb2da5",
   656 => x"a45188eb",
   657 => x"2da4b851",
   658 => x"88eb2da7",
   659 => x"8408a5e4",
   660 => x"08705471",
   661 => x"87e82953",
   662 => x"5b569a87",
   663 => x"2d8808a6",
   664 => x"fc0c7552",
   665 => x"7987e829",
   666 => x"519a872d",
   667 => x"8808a780",
   668 => x"0c755279",
   669 => x"84b92951",
   670 => x"9a872d88",
   671 => x"0880f6b4",
   672 => x"0ca3b451",
   673 => x"88eb2da6",
   674 => x"fc0852a3",
   675 => x"e45188eb",
   676 => x"2da3ec51",
   677 => x"88eb2da7",
   678 => x"800852a3",
   679 => x"e45188eb",
   680 => x"2d80f6b4",
   681 => x"0852a49c",
   682 => x"5188eb2d",
   683 => x"a4b85188",
   684 => x"eb2d800b",
   685 => x"880c02b8",
   686 => x"050d0402",
   687 => x"b805f805",
   688 => x"52805196",
   689 => x"ad2d9f53",
   690 => x"a5c45280",
   691 => x"f690519e",
   692 => x"e52d7778",
   693 => x"80f6840c",
   694 => x"81177081",
   695 => x"ff0680f6",
   696 => x"8c0b84e0",
   697 => x"2d525856",
   698 => x"5a92ea04",
   699 => x"760856b0",
   700 => x"53755276",
   701 => x"519ee52d",
   702 => x"80c10b80",
   703 => x"f68c0b84",
   704 => x"e02d5656",
   705 => x"92c604ff",
   706 => x"15707831",
   707 => x"7c0c5980",
   708 => x"59939704",
   709 => x"02f8050d",
   710 => x"73823270",
   711 => x"09810570",
   712 => x"72078025",
   713 => x"880c5252",
   714 => x"0288050d",
   715 => x"0402f405",
   716 => x"0d747671",
   717 => x"53545271",
   718 => x"822e8338",
   719 => x"83517181",
   720 => x"2e9b3881",
   721 => x"7226a038",
   722 => x"71822ebc",
   723 => x"3871842e",
   724 => x"ac387073",
   725 => x"0c70880c",
   726 => x"028c050d",
   727 => x"0480e40b",
   728 => x"80f68408",
   729 => x"258c3880",
   730 => x"730c7088",
   731 => x"0c028c05",
   732 => x"0d048373",
   733 => x"0c70880c",
   734 => x"028c050d",
   735 => x"0482730c",
   736 => x"70880c02",
   737 => x"8c050d04",
   738 => x"81730c70",
   739 => x"880c028c",
   740 => x"050d0402",
   741 => x"fc050d74",
   742 => x"74148205",
   743 => x"710c880c",
   744 => x"0284050d",
   745 => x"0402d805",
   746 => x"0d7b7d7f",
   747 => x"61851270",
   748 => x"822b7511",
   749 => x"70747170",
   750 => x"8405530c",
   751 => x"5a5a5d5b",
   752 => x"760c7980",
   753 => x"f8180c79",
   754 => x"86125257",
   755 => x"585a5a76",
   756 => x"76249938",
   757 => x"76b32982",
   758 => x"2b791151",
   759 => x"53767370",
   760 => x"8405550c",
   761 => x"81145475",
   762 => x"7425f238",
   763 => x"7681cc29",
   764 => x"19fc1108",
   765 => x"8105fc12",
   766 => x"0c7a1970",
   767 => x"089fa013",
   768 => x"0c585685",
   769 => x"0b80f684",
   770 => x"0c75880c",
   771 => x"02a8050d",
   772 => x"0402f405",
   773 => x"0d029305",
   774 => x"84e02d51",
   775 => x"80028405",
   776 => x"970584e0",
   777 => x"2d545270",
   778 => x"732e8938",
   779 => x"71880c02",
   780 => x"8c050d04",
   781 => x"7080f688",
   782 => x"0b85802d",
   783 => x"810b880c",
   784 => x"028c050d",
   785 => x"0402dc05",
   786 => x"0d7a7c59",
   787 => x"56820b83",
   788 => x"19555574",
   789 => x"167084e0",
   790 => x"2d7584e0",
   791 => x"2d5b5153",
   792 => x"72792e80",
   793 => x"c73880c1",
   794 => x"0b811681",
   795 => x"16565657",
   796 => x"827525df",
   797 => x"38ffa917",
   798 => x"7081ff06",
   799 => x"55597382",
   800 => x"26833887",
   801 => x"55815376",
   802 => x"80d22e98",
   803 => x"38775275",
   804 => x"519ffe2d",
   805 => x"80537288",
   806 => x"08258938",
   807 => x"871580f6",
   808 => x"840c8153",
   809 => x"72880c02",
   810 => x"a4050d04",
   811 => x"7280f688",
   812 => x"0b85802d",
   813 => x"827525ff",
   814 => x"9a3898f5",
   815 => x"04940802",
   816 => x"940cfd3d",
   817 => x"0d805394",
   818 => x"088c0508",
   819 => x"52940888",
   820 => x"05085182",
   821 => x"de3f8808",
   822 => x"70880c54",
   823 => x"853d0d94",
   824 => x"0c049408",
   825 => x"02940cfd",
   826 => x"3d0d8153",
   827 => x"94088c05",
   828 => x"08529408",
   829 => x"88050851",
   830 => x"82b93f88",
   831 => x"0870880c",
   832 => x"54853d0d",
   833 => x"940c0494",
   834 => x"0802940c",
   835 => x"f93d0d80",
   836 => x"0b9408fc",
   837 => x"050c9408",
   838 => x"88050880",
   839 => x"25ab3894",
   840 => x"08880508",
   841 => x"30940888",
   842 => x"050c800b",
   843 => x"9408f405",
   844 => x"0c9408fc",
   845 => x"05088838",
   846 => x"810b9408",
   847 => x"f4050c94",
   848 => x"08f40508",
   849 => x"9408fc05",
   850 => x"0c94088c",
   851 => x"05088025",
   852 => x"ab389408",
   853 => x"8c050830",
   854 => x"94088c05",
   855 => x"0c800b94",
   856 => x"08f0050c",
   857 => x"9408fc05",
   858 => x"08883881",
   859 => x"0b9408f0",
   860 => x"050c9408",
   861 => x"f0050894",
   862 => x"08fc050c",
   863 => x"80539408",
   864 => x"8c050852",
   865 => x"94088805",
   866 => x"085181a7",
   867 => x"3f880870",
   868 => x"9408f805",
   869 => x"0c549408",
   870 => x"fc050880",
   871 => x"2e8c3894",
   872 => x"08f80508",
   873 => x"309408f8",
   874 => x"050c9408",
   875 => x"f8050870",
   876 => x"880c5489",
   877 => x"3d0d940c",
   878 => x"04940802",
   879 => x"940cfb3d",
   880 => x"0d800b94",
   881 => x"08fc050c",
   882 => x"94088805",
   883 => x"08802593",
   884 => x"38940888",
   885 => x"05083094",
   886 => x"0888050c",
   887 => x"810b9408",
   888 => x"fc050c94",
   889 => x"088c0508",
   890 => x"80258c38",
   891 => x"94088c05",
   892 => x"08309408",
   893 => x"8c050c81",
   894 => x"5394088c",
   895 => x"05085294",
   896 => x"08880508",
   897 => x"51ad3f88",
   898 => x"08709408",
   899 => x"f8050c54",
   900 => x"9408fc05",
   901 => x"08802e8c",
   902 => x"389408f8",
   903 => x"05083094",
   904 => x"08f8050c",
   905 => x"9408f805",
   906 => x"0870880c",
   907 => x"54873d0d",
   908 => x"940c0494",
   909 => x"0802940c",
   910 => x"fd3d0d81",
   911 => x"0b9408fc",
   912 => x"050c800b",
   913 => x"9408f805",
   914 => x"0c94088c",
   915 => x"05089408",
   916 => x"88050827",
   917 => x"ac389408",
   918 => x"fc050880",
   919 => x"2ea33880",
   920 => x"0b94088c",
   921 => x"05082499",
   922 => x"3894088c",
   923 => x"05081094",
   924 => x"088c050c",
   925 => x"9408fc05",
   926 => x"08109408",
   927 => x"fc050cc9",
   928 => x"399408fc",
   929 => x"0508802e",
   930 => x"80c93894",
   931 => x"088c0508",
   932 => x"94088805",
   933 => x"0826a138",
   934 => x"94088805",
   935 => x"0894088c",
   936 => x"05083194",
   937 => x"0888050c",
   938 => x"9408f805",
   939 => x"089408fc",
   940 => x"05080794",
   941 => x"08f8050c",
   942 => x"9408fc05",
   943 => x"08812a94",
   944 => x"08fc050c",
   945 => x"94088c05",
   946 => x"08812a94",
   947 => x"088c050c",
   948 => x"ffaf3994",
   949 => x"08900508",
   950 => x"802e8f38",
   951 => x"94088805",
   952 => x"08709408",
   953 => x"f4050c51",
   954 => x"8d399408",
   955 => x"f8050870",
   956 => x"9408f405",
   957 => x"0c519408",
   958 => x"f4050888",
   959 => x"0c853d0d",
   960 => x"940c0494",
   961 => x"0802940c",
   962 => x"ff3d0d80",
   963 => x"0b9408fc",
   964 => x"050c9408",
   965 => x"88050881",
   966 => x"06ff1170",
   967 => x"09709408",
   968 => x"8c050806",
   969 => x"9408fc05",
   970 => x"08119408",
   971 => x"fc050c94",
   972 => x"08880508",
   973 => x"812a9408",
   974 => x"88050c94",
   975 => x"088c0508",
   976 => x"1094088c",
   977 => x"050c5151",
   978 => x"51519408",
   979 => x"88050880",
   980 => x"2e8438ff",
   981 => x"bd399408",
   982 => x"fc050870",
   983 => x"880c5183",
   984 => x"3d0d940c",
   985 => x"04fc3d0d",
   986 => x"7670797b",
   987 => x"55555555",
   988 => x"8f72278c",
   989 => x"38727507",
   990 => x"83065170",
   991 => x"802ea738",
   992 => x"ff125271",
   993 => x"ff2e9838",
   994 => x"72708105",
   995 => x"54337470",
   996 => x"81055634",
   997 => x"ff125271",
   998 => x"ff2e0981",
   999 => x"06ea3874",
  1000 => x"880c863d",
  1001 => x"0d047451",
  1002 => x"72708405",
  1003 => x"54087170",
  1004 => x"8405530c",
  1005 => x"72708405",
  1006 => x"54087170",
  1007 => x"8405530c",
  1008 => x"72708405",
  1009 => x"54087170",
  1010 => x"8405530c",
  1011 => x"72708405",
  1012 => x"54087170",
  1013 => x"8405530c",
  1014 => x"f0125271",
  1015 => x"8f26c938",
  1016 => x"83722795",
  1017 => x"38727084",
  1018 => x"05540871",
  1019 => x"70840553",
  1020 => x"0cfc1252",
  1021 => x"718326ed",
  1022 => x"387054ff",
  1023 => x"8339fb3d",
  1024 => x"0d777970",
  1025 => x"72078306",
  1026 => x"53545270",
  1027 => x"93387173",
  1028 => x"73085456",
  1029 => x"54717308",
  1030 => x"2e80c438",
  1031 => x"73755452",
  1032 => x"71337081",
  1033 => x"ff065254",
  1034 => x"70802e9d",
  1035 => x"38723355",
  1036 => x"70752e09",
  1037 => x"81069538",
  1038 => x"81128114",
  1039 => x"71337081",
  1040 => x"ff065456",
  1041 => x"545270e5",
  1042 => x"38723355",
  1043 => x"7381ff06",
  1044 => x"7581ff06",
  1045 => x"71713188",
  1046 => x"0c525287",
  1047 => x"3d0d0471",
  1048 => x"0970f7fb",
  1049 => x"fdff1406",
  1050 => x"70f88482",
  1051 => x"81800651",
  1052 => x"51517097",
  1053 => x"38841484",
  1054 => x"16710854",
  1055 => x"56547175",
  1056 => x"082edc38",
  1057 => x"73755452",
  1058 => x"ff963980",
  1059 => x"0b880c87",
  1060 => x"3d0d0400",
  1061 => x"00ffffff",
  1062 => x"ff00ffff",
  1063 => x"ffff00ff",
  1064 => x"ffffff00",
  1065 => x"30313233",
  1066 => x"34353637",
  1067 => x"38394142",
  1068 => x"43444546",
  1069 => x"00000000",
  1070 => x"44485259",
  1071 => x"53544f4e",
  1072 => x"45205052",
  1073 => x"4f475241",
  1074 => x"4d2c2053",
  1075 => x"4f4d4520",
  1076 => x"53545249",
  1077 => x"4e470000",
  1078 => x"44485259",
  1079 => x"53544f4e",
  1080 => x"45205052",
  1081 => x"4f475241",
  1082 => x"4d2c2031",
  1083 => x"27535420",
  1084 => x"53545249",
  1085 => x"4e470000",
  1086 => x"44687279",
  1087 => x"73746f6e",
  1088 => x"65204265",
  1089 => x"6e63686d",
  1090 => x"61726b2c",
  1091 => x"20566572",
  1092 => x"73696f6e",
  1093 => x"20322e31",
  1094 => x"20284c61",
  1095 => x"6e677561",
  1096 => x"67653a20",
  1097 => x"43290a00",
  1098 => x"50726f67",
  1099 => x"72616d20",
  1100 => x"636f6d70",
  1101 => x"696c6564",
  1102 => x"20776974",
  1103 => x"68202772",
  1104 => x"65676973",
  1105 => x"74657227",
  1106 => x"20617474",
  1107 => x"72696275",
  1108 => x"74650a00",
  1109 => x"45786563",
  1110 => x"7574696f",
  1111 => x"6e207374",
  1112 => x"61727473",
  1113 => x"2c202564",
  1114 => x"2072756e",
  1115 => x"73207468",
  1116 => x"726f7567",
  1117 => x"68204468",
  1118 => x"72797374",
  1119 => x"6f6e650a",
  1120 => x"00000000",
  1121 => x"44485259",
  1122 => x"53544f4e",
  1123 => x"45205052",
  1124 => x"4f475241",
  1125 => x"4d2c2032",
  1126 => x"274e4420",
  1127 => x"53545249",
  1128 => x"4e470000",
  1129 => x"55736572",
  1130 => x"2074696d",
  1131 => x"653a2025",
  1132 => x"640a0000",
  1133 => x"4d696372",
  1134 => x"6f736563",
  1135 => x"6f6e6473",
  1136 => x"20666f72",
  1137 => x"206f6e65",
  1138 => x"2072756e",
  1139 => x"20746872",
  1140 => x"6f756768",
  1141 => x"20446872",
  1142 => x"7973746f",
  1143 => x"6e653a20",
  1144 => x"00000000",
  1145 => x"2564200a",
  1146 => x"00000000",
  1147 => x"44687279",
  1148 => x"73746f6e",
  1149 => x"65732070",
  1150 => x"65722053",
  1151 => x"65636f6e",
  1152 => x"643a2020",
  1153 => x"20202020",
  1154 => x"20202020",
  1155 => x"20202020",
  1156 => x"20202020",
  1157 => x"20202020",
  1158 => x"00000000",
  1159 => x"56415820",
  1160 => x"4d495053",
  1161 => x"20726174",
  1162 => x"696e6720",
  1163 => x"2a203130",
  1164 => x"3030203d",
  1165 => x"20256420",
  1166 => x"0a000000",
  1167 => x"50726f67",
  1168 => x"72616d20",
  1169 => x"636f6d70",
  1170 => x"696c6564",
  1171 => x"20776974",
  1172 => x"686f7574",
  1173 => x"20277265",
  1174 => x"67697374",
  1175 => x"65722720",
  1176 => x"61747472",
  1177 => x"69627574",
  1178 => x"650a0000",
  1179 => x"4d656173",
  1180 => x"75726564",
  1181 => x"2074696d",
  1182 => x"6520746f",
  1183 => x"6f20736d",
  1184 => x"616c6c20",
  1185 => x"746f206f",
  1186 => x"62746169",
  1187 => x"6e206d65",
  1188 => x"616e696e",
  1189 => x"6766756c",
  1190 => x"20726573",
  1191 => x"756c7473",
  1192 => x"0a000000",
  1193 => x"506c6561",
  1194 => x"73652069",
  1195 => x"6e637265",
  1196 => x"61736520",
  1197 => x"6e756d62",
  1198 => x"6572206f",
  1199 => x"66207275",
  1200 => x"6e730a00",
  1201 => x"44485259",
  1202 => x"53544f4e",
  1203 => x"45205052",
  1204 => x"4f475241",
  1205 => x"4d2c2033",
  1206 => x"27524420",
  1207 => x"53545249",
  1208 => x"4e470000",
  1209 => x"000061a8",
  1210 => x"00000000",
	others => x"00000000"
);

begin

process (clk)
begin
	if (clk'event and clk = '1') then
		if (from_zpu.memAWriteEnable = '1') and (from_zpu.memBWriteEnable = '1') and (from_zpu.memAAddr=from_zpu.memBAddr) and (from_zpu.memAWrite/=from_zpu.memBWrite) then
			report "write collision" severity failure;
		end if;
	
		if (from_zpu.memAWriteEnable = '1') then
			ram(to_integer(unsigned(from_zpu.memAAddr(maxAddrBit downto 2)))) := from_zpu.memAWrite;
			to_zpu.memARead <= from_zpu.memAWrite;
		else
			to_zpu.memARead <= ram(to_integer(unsigned(from_zpu.memAAddr(maxAddrBit downto 2))));
		end if;
	end if;
end process;

process (clk)
begin
	if (clk'event and clk = '1') then
		if (from_zpu.memBWriteEnable = '1') then
			ram(to_integer(unsigned(from_zpu.memBAddr(maxAddrBit downto 2)))) := from_zpu.memBWrite;
			to_zpu.memBRead <= from_zpu.memBWrite;
		else
			to_zpu.memBRead <= ram(to_integer(unsigned(from_zpu.memBAddr(maxAddrBit downto 2))));
		end if;
	end if;
end process;


end arch;

