-- ZPU
--
-- Copyright 2004-2008 oharboe - �yvind Harboe - oyvind.harboe@zylin.com
-- Modified by Alastair M. Robinson for the ZPUFlex project.
--
-- The FreeBSD license
-- 
-- Redistribution and use in source and binary forms, with or without
-- modification, are permitted provided that the following conditions
-- are met:
-- 
-- 1. Redistributions of source code must retain the above copyright
--    notice, this list of conditions and the following disclaimer.
-- 2. Redistributions in binary form must reproduce the above
--    copyright notice, this list of conditions and the following
--    disclaimer in the documentation and/or other materials
--    provided with the distribution.
-- 
-- THIS SOFTWARE IS PROVIDED BY THE ZPU PROJECT ``AS IS'' AND ANY
-- EXPRESS OR IMPLIED WARRANTIES, INCLUDING, BUT NOT LIMITED TO,
-- THE IMPLIED WARRANTIES OF MERCHANTABILITY AND FITNESS FOR A
-- PARTICULAR PURPOSE ARE DISCLAIMED. IN NO EVENT SHALL THE
-- ZPU PROJECT OR CONTRIBUTORS BE LIABLE FOR ANY DIRECT,
-- INDIRECT, INCIDENTAL, SPECIAL, EXEMPLARY, OR CONSEQUENTIAL DAMAGES
-- (INCLUDING, BUT NOT LIMITED TO, PROCUREMENT OF SUBSTITUTE GOODS
-- OR SERVICES; LOSS OF USE, DATA, OR PROFITS; OR BUSINESS INTERRUPTION)
-- HOWEVER CAUSED AND ON ANY THEORY OF LIABILITY, WHETHER IN CONTRACT,
-- STRICT LIABILITY, OR TORT (INCLUDING NEGLIGENCE OR OTHERWISE)
-- ARISING IN ANY WAY OUT OF THE USE OF THIS SOFTWARE, EVEN IF
-- ADVISED OF THE POSSIBILITY OF SUCH DAMAGE.
-- 
-- The views and conclusions contained in the software and documentation
-- are those of the authors and should not be interpreted as representing
-- official policies, either expressed or implied, of the ZPU Project.

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;


library work;
use work.zpupkg.all;

entity VGATest_ROM is
generic
	(
		maxAddrBitBRAM : integer := maxAddrBitBRAMLimit -- Specify your actual ROM size to save LEs and unnecessary block RAM usage.
	);
port (
	clk : in std_logic;
	areset : in std_logic := '0';
	from_zpu : in ZPU_ToROM;
	to_zpu : out ZPU_FromROM
);
end VGATest_ROM;

architecture arch of VGATest_ROM is

type ram_type is array(natural range 0 to ((2**(maxAddrBitBRAM+1))/4)-1) of std_logic_vector(wordSize-1 downto 0);

shared variable ram : ram_type :=
(
     0 => x"84808080",
     1 => x"ee040000",
     2 => x"00000000",
     3 => x"84808080",
     4 => x"88080d80",
     5 => x"04848080",
     6 => x"80950471",
     7 => x"fd060872",
     8 => x"83060981",
     9 => x"05820583",
    10 => x"2b2a83ff",
    11 => x"ff065204",
    12 => x"71fc0608",
    13 => x"72830609",
    14 => x"81058305",
    15 => x"1010102a",
    16 => x"81ff0652",
    17 => x"0471fc06",
    18 => x"08848080",
    19 => x"92c47383",
    20 => x"06101005",
    21 => x"08067381",
    22 => x"ff067383",
    23 => x"06098105",
    24 => x"83051010",
    25 => x"102b0772",
    26 => x"fc060c51",
    27 => x"51040284",
    28 => x"05848080",
    29 => x"80880c84",
    30 => x"80808095",
    31 => x"0b848080",
    32 => x"85f80400",
    33 => x"02c0050d",
    34 => x"0280c405",
    35 => x"5b80707c",
    36 => x"7084055e",
    37 => x"08725f5f",
    38 => x"5f5a7c70",
    39 => x"84055e08",
    40 => x"57805976",
    41 => x"982a7788",
    42 => x"2b585574",
    43 => x"802e82f3",
    44 => x"387b802e",
    45 => x"80d33880",
    46 => x"5c7480e4",
    47 => x"2e81de38",
    48 => x"7480f82e",
    49 => x"81d73874",
    50 => x"80e42e81",
    51 => x"e2387480",
    52 => x"e42680f1",
    53 => x"387480e3",
    54 => x"2e80c838",
    55 => x"a5518480",
    56 => x"8085882d",
    57 => x"74518480",
    58 => x"8085882d",
    59 => x"821a811a",
    60 => x"5a5a8379",
    61 => x"25ffac38",
    62 => x"74ff9f38",
    63 => x"7e848080",
    64 => x"98d00c02",
    65 => x"80c0050d",
    66 => x"0474a52e",
    67 => x"0981069b",
    68 => x"38810b81",
    69 => x"1a5a5c83",
    70 => x"7925ff87",
    71 => x"38848080",
    72 => x"81f8047a",
    73 => x"841c7108",
    74 => x"575c5474",
    75 => x"51848080",
    76 => x"85882d81",
    77 => x"1a811a5a",
    78 => x"5a837925",
    79 => x"fee53884",
    80 => x"808081f8",
    81 => x"047480f3",
    82 => x"2e81e538",
    83 => x"7480f82e",
    84 => x"098106ff",
    85 => x"87387d53",
    86 => x"8058777e",
    87 => x"24829638",
    88 => x"72802e81",
    89 => x"f9388756",
    90 => x"729c2a73",
    91 => x"842b5452",
    92 => x"71802e83",
    93 => x"388158b7",
    94 => x"12547189",
    95 => x"248438b0",
    96 => x"12547780",
    97 => x"f038ff16",
    98 => x"56758025",
    99 => x"db388119",
   100 => x"59837925",
   101 => x"fe8d3884",
   102 => x"808081f8",
   103 => x"047a841c",
   104 => x"7108405c",
   105 => x"527480e4",
   106 => x"2e098106",
   107 => x"fea0387d",
   108 => x"54805877",
   109 => x"7e248195",
   110 => x"3873802e",
   111 => x"81a03887",
   112 => x"56739c2a",
   113 => x"74842b55",
   114 => x"5271802e",
   115 => x"83388158",
   116 => x"b7125371",
   117 => x"89248438",
   118 => x"b0125377",
   119 => x"af38ff16",
   120 => x"56758025",
   121 => x"dc388119",
   122 => x"59837925",
   123 => x"fdb53884",
   124 => x"808081f8",
   125 => x"04735184",
   126 => x"80808588",
   127 => x"2dff1656",
   128 => x"758025fe",
   129 => x"e3388480",
   130 => x"80838e04",
   131 => x"72518480",
   132 => x"8085882d",
   133 => x"ff165675",
   134 => x"8025ffa5",
   135 => x"38848080",
   136 => x"83e60479",
   137 => x"84808098",
   138 => x"d00c0280",
   139 => x"c0050d04",
   140 => x"7a841c71",
   141 => x"08535c53",
   142 => x"84808085",
   143 => x"ad2d8119",
   144 => x"59837925",
   145 => x"fcdd3884",
   146 => x"808081f8",
   147 => x"04ad5184",
   148 => x"80808588",
   149 => x"2d7d0981",
   150 => x"055473fe",
   151 => x"e238b051",
   152 => x"84808085",
   153 => x"882d8119",
   154 => x"59837925",
   155 => x"fcb53884",
   156 => x"808081f8",
   157 => x"04ad5184",
   158 => x"80808588",
   159 => x"2d7d0981",
   160 => x"05538480",
   161 => x"8082e004",
   162 => x"02f8050d",
   163 => x"7352c008",
   164 => x"70882a70",
   165 => x"81065151",
   166 => x"5170802e",
   167 => x"f13871c0",
   168 => x"0c718480",
   169 => x"8098d00c",
   170 => x"0288050d",
   171 => x"0402e805",
   172 => x"0d807857",
   173 => x"55757084",
   174 => x"05570853",
   175 => x"80547298",
   176 => x"2a73882b",
   177 => x"54527180",
   178 => x"2ea238c0",
   179 => x"0870882a",
   180 => x"70810651",
   181 => x"51517080",
   182 => x"2ef13871",
   183 => x"c00c8115",
   184 => x"81155555",
   185 => x"837425d6",
   186 => x"3871ca38",
   187 => x"74848080",
   188 => x"98d00c02",
   189 => x"98050d04",
   190 => x"02dc050d",
   191 => x"80528480",
   192 => x"800bfc80",
   193 => x"0c811270",
   194 => x"55598480",
   195 => x"80568055",
   196 => x"84fe5381",
   197 => x"1483ffff",
   198 => x"06707770",
   199 => x"8405590c",
   200 => x"fe145454",
   201 => x"728025eb",
   202 => x"38811555",
   203 => x"83df7525",
   204 => x"df388057",
   205 => x"805584fe",
   206 => x"53fc8008",
   207 => x"fe145452",
   208 => x"728025f5",
   209 => x"38811555",
   210 => x"83df7525",
   211 => x"e9388117",
   212 => x"57b17725",
   213 => x"df388058",
   214 => x"75558057",
   215 => x"84fe5381",
   216 => x"1483ffff",
   217 => x"06707670",
   218 => x"8405580c",
   219 => x"fe145454",
   220 => x"728025eb",
   221 => x"38811757",
   222 => x"83df7725",
   223 => x"df388118",
   224 => x"58937825",
   225 => x"d3388119",
   226 => x"52805184",
   227 => x"80808f81",
   228 => x"2d848080",
   229 => x"86850402",
   230 => x"f4050d74",
   231 => x"76525380",
   232 => x"71259038",
   233 => x"70527270",
   234 => x"84055408",
   235 => x"ff135351",
   236 => x"71f43802",
   237 => x"8c050d04",
   238 => x"02d4050d",
   239 => x"7c7e5c58",
   240 => x"810b8480",
   241 => x"8092d458",
   242 => x"5a835976",
   243 => x"08780c77",
   244 => x"08770856",
   245 => x"5473752e",
   246 => x"94387708",
   247 => x"53745284",
   248 => x"808092e4",
   249 => x"51848080",
   250 => x"81842d80",
   251 => x"5a775680",
   252 => x"7b259038",
   253 => x"7a557570",
   254 => x"84055708",
   255 => x"ff165654",
   256 => x"74f43877",
   257 => x"08770856",
   258 => x"5675752e",
   259 => x"94387708",
   260 => x"53745284",
   261 => x"808093a4",
   262 => x"51848080",
   263 => x"81842d80",
   264 => x"5aff1984",
   265 => x"18585978",
   266 => x"8025ff9f",
   267 => x"38798480",
   268 => x"8098d00c",
   269 => x"02ac050d",
   270 => x"0402e405",
   271 => x"0d787a55",
   272 => x"56815785",
   273 => x"aad5aad5",
   274 => x"760cfad5",
   275 => x"aad5aa0b",
   276 => x"8c170ccc",
   277 => x"76848080",
   278 => x"80c52db3",
   279 => x"0b8f1784",
   280 => x"808080c5",
   281 => x"2d750853",
   282 => x"72fce2d5",
   283 => x"aad52e92",
   284 => x"38750852",
   285 => x"84808093",
   286 => x"e4518480",
   287 => x"8081842d",
   288 => x"80578c16",
   289 => x"085574fa",
   290 => x"d5aad4b3",
   291 => x"2e93388c",
   292 => x"16085284",
   293 => x"808094a0",
   294 => x"51848080",
   295 => x"81842d80",
   296 => x"57755580",
   297 => x"74258e38",
   298 => x"74708405",
   299 => x"5608ff15",
   300 => x"555373f4",
   301 => x"38750854",
   302 => x"73fce2d5",
   303 => x"aad52e92",
   304 => x"38750852",
   305 => x"84808094",
   306 => x"dc518480",
   307 => x"8081842d",
   308 => x"80578c16",
   309 => x"085372fa",
   310 => x"d5aad4b3",
   311 => x"2e93388c",
   312 => x"16085284",
   313 => x"80809598",
   314 => x"51848080",
   315 => x"81842d80",
   316 => x"57768480",
   317 => x"8098d00c",
   318 => x"029c050d",
   319 => x"0402c405",
   320 => x"0d605b80",
   321 => x"62908080",
   322 => x"29ff0584",
   323 => x"808095d4",
   324 => x"53405a84",
   325 => x"80808184",
   326 => x"2d80e1b3",
   327 => x"5780fe5e",
   328 => x"ae518480",
   329 => x"8085882d",
   330 => x"76107096",
   331 => x"2a810656",
   332 => x"5774802e",
   333 => x"85387681",
   334 => x"07577695",
   335 => x"2a810658",
   336 => x"77802e85",
   337 => x"38768132",
   338 => x"57787707",
   339 => x"7f06775e",
   340 => x"598fffff",
   341 => x"5876bfff",
   342 => x"ff06707a",
   343 => x"32822b7c",
   344 => x"11515776",
   345 => x"0c761070",
   346 => x"962a8106",
   347 => x"56577480",
   348 => x"2e853876",
   349 => x"81075776",
   350 => x"952a8106",
   351 => x"5574802e",
   352 => x"85387681",
   353 => x"3257ff18",
   354 => x"58778025",
   355 => x"c8387c57",
   356 => x"8fffff58",
   357 => x"76bfffff",
   358 => x"06707a32",
   359 => x"822b7c05",
   360 => x"7008575e",
   361 => x"5674762e",
   362 => x"80ea3880",
   363 => x"7a538480",
   364 => x"8095e452",
   365 => x"5c848080",
   366 => x"81842d74",
   367 => x"54755375",
   368 => x"52848080",
   369 => x"95f85184",
   370 => x"80808184",
   371 => x"2d7b5a76",
   372 => x"1070962a",
   373 => x"81065757",
   374 => x"75802e85",
   375 => x"38768107",
   376 => x"5776952a",
   377 => x"81065574",
   378 => x"802e8538",
   379 => x"76813257",
   380 => x"ff185877",
   381 => x"8025ff9c",
   382 => x"38ff1e5e",
   383 => x"7dfea138",
   384 => x"8a518480",
   385 => x"8085882d",
   386 => x"7b848080",
   387 => x"98d00c02",
   388 => x"bc050d04",
   389 => x"811a5a84",
   390 => x"80808bcf",
   391 => x"0402cc05",
   392 => x"0d7e605e",
   393 => x"58815a80",
   394 => x"5b80c07a",
   395 => x"585c85ad",
   396 => x"a989bb78",
   397 => x"0c795981",
   398 => x"56975576",
   399 => x"7607822b",
   400 => x"78115154",
   401 => x"85ada989",
   402 => x"bb740c75",
   403 => x"10ff1656",
   404 => x"56748025",
   405 => x"e6387610",
   406 => x"811a5a57",
   407 => x"987925d7",
   408 => x"38775680",
   409 => x"7d259038",
   410 => x"7c557570",
   411 => x"84055708",
   412 => x"ff165654",
   413 => x"74f43881",
   414 => x"57ff8787",
   415 => x"a5c3780c",
   416 => x"97597682",
   417 => x"2b781170",
   418 => x"085f5656",
   419 => x"7cff8787",
   420 => x"a5c32e80",
   421 => x"cc387408",
   422 => x"547385ad",
   423 => x"a989bb2e",
   424 => x"94388075",
   425 => x"08547653",
   426 => x"84808096",
   427 => x"a0525a84",
   428 => x"80808184",
   429 => x"2d7610ff",
   430 => x"1a5a5778",
   431 => x"8025c338",
   432 => x"7a822b56",
   433 => x"75b1387b",
   434 => x"52848080",
   435 => x"96c05184",
   436 => x"80808184",
   437 => x"2d7b8480",
   438 => x"8098d00c",
   439 => x"02b4050d",
   440 => x"047a7707",
   441 => x"7710ff1b",
   442 => x"5b585b78",
   443 => x"8025ff92",
   444 => x"38848080",
   445 => x"8dc00475",
   446 => x"52848080",
   447 => x"96fc5184",
   448 => x"80808184",
   449 => x"2d75992a",
   450 => x"81328106",
   451 => x"70098105",
   452 => x"71077009",
   453 => x"709f2c7d",
   454 => x"0679109f",
   455 => x"fffffc06",
   456 => x"60812a41",
   457 => x"5a5d5758",
   458 => x"5975da38",
   459 => x"79098105",
   460 => x"707b079f",
   461 => x"2a55567b",
   462 => x"bf268438",
   463 => x"739d3881",
   464 => x"70538480",
   465 => x"8096c052",
   466 => x"5c848080",
   467 => x"81842d7b",
   468 => x"84808098",
   469 => x"d00c02b4",
   470 => x"050d0484",
   471 => x"80809794",
   472 => x"51848080",
   473 => x"81842d7b",
   474 => x"52848080",
   475 => x"96c05184",
   476 => x"80808184",
   477 => x"2d7b8480",
   478 => x"8098d00c",
   479 => x"02b4050d",
   480 => x"0402d405",
   481 => x"0d7c5781",
   482 => x"70848080",
   483 => x"92d45b59",
   484 => x"5b835a78",
   485 => x"08770c76",
   486 => x"08790856",
   487 => x"5473752e",
   488 => x"94387608",
   489 => x"53745284",
   490 => x"808092e4",
   491 => x"51848080",
   492 => x"81842d80",
   493 => x"5876569f",
   494 => x"ff557570",
   495 => x"84055708",
   496 => x"ff165654",
   497 => x"748025f2",
   498 => x"38760879",
   499 => x"08565675",
   500 => x"752e9438",
   501 => x"76085374",
   502 => x"52848080",
   503 => x"93a45184",
   504 => x"80808184",
   505 => x"2d8058ff",
   506 => x"1a841a5a",
   507 => x"5a798025",
   508 => x"ffa13877",
   509 => x"81fd3877",
   510 => x"5b815885",
   511 => x"aad5aad5",
   512 => x"770cfad5",
   513 => x"aad5aa0b",
   514 => x"8c180ccc",
   515 => x"77848080",
   516 => x"80c52db3",
   517 => x"0b8f1884",
   518 => x"808080c5",
   519 => x"2d760855",
   520 => x"74fce2d5",
   521 => x"aad52e92",
   522 => x"38760852",
   523 => x"84808093",
   524 => x"e4518480",
   525 => x"8081842d",
   526 => x"80588c17",
   527 => x"085978fa",
   528 => x"d5aad4b3",
   529 => x"2e93388c",
   530 => x"17085284",
   531 => x"808094a0",
   532 => x"51848080",
   533 => x"81842d80",
   534 => x"5876569f",
   535 => x"ff557570",
   536 => x"84055708",
   537 => x"ff165654",
   538 => x"748025f2",
   539 => x"3876085a",
   540 => x"79fce2d5",
   541 => x"aad52e92",
   542 => x"38760852",
   543 => x"84808094",
   544 => x"dc518480",
   545 => x"8081842d",
   546 => x"80588c17",
   547 => x"085473fa",
   548 => x"d5aad4b3",
   549 => x"2e80ee38",
   550 => x"8c170852",
   551 => x"84808095",
   552 => x"98518480",
   553 => x"8081842d",
   554 => x"8058775b",
   555 => x"a0805276",
   556 => x"51848080",
   557 => x"8c9d2d84",
   558 => x"808098d0",
   559 => x"08548480",
   560 => x"8098d008",
   561 => x"80e93884",
   562 => x"808098d0",
   563 => x"085b7352",
   564 => x"76518480",
   565 => x"8089fd2d",
   566 => x"84808098",
   567 => x"d008be38",
   568 => x"84808098",
   569 => x"d0085b7a",
   570 => x"84808098",
   571 => x"d00c02ac",
   572 => x"050d0484",
   573 => x"808097e0",
   574 => x"51848080",
   575 => x"81842d84",
   576 => x"80808ff9",
   577 => x"0477802e",
   578 => x"ffa03884",
   579 => x"80809884",
   580 => x"51848080",
   581 => x"81842d84",
   582 => x"808091ac",
   583 => x"04848080",
   584 => x"98a05184",
   585 => x"80808184",
   586 => x"2d848080",
   587 => x"91e70484",
   588 => x"808098b8",
   589 => x"51848080",
   590 => x"81842d84",
   591 => x"808091ce",
   592 => x"04000000",
   593 => x"00ffffff",
   594 => x"ff00ffff",
   595 => x"ffff00ff",
   596 => x"ffffff00",
   597 => x"00000000",
   598 => x"55555555",
   599 => x"aaaaaaaa",
   600 => x"ffffffff",
   601 => x"53616e69",
   602 => x"74792063",
   603 => x"6865636b",
   604 => x"20666169",
   605 => x"6c656420",
   606 => x"28626566",
   607 => x"6f726520",
   608 => x"63616368",
   609 => x"65207265",
   610 => x"66726573",
   611 => x"6829206f",
   612 => x"6e203078",
   613 => x"25642028",
   614 => x"676f7420",
   615 => x"30782564",
   616 => x"290a0000",
   617 => x"53616e69",
   618 => x"74792063",
   619 => x"6865636b",
   620 => x"20666169",
   621 => x"6c656420",
   622 => x"28616674",
   623 => x"65722063",
   624 => x"61636865",
   625 => x"20726566",
   626 => x"72657368",
   627 => x"29206f6e",
   628 => x"20307825",
   629 => x"64202867",
   630 => x"6f742030",
   631 => x"78256429",
   632 => x"0a000000",
   633 => x"42797465",
   634 => x"20636865",
   635 => x"636b2066",
   636 => x"61696c65",
   637 => x"64202862",
   638 => x"65666f72",
   639 => x"65206361",
   640 => x"63686520",
   641 => x"72656672",
   642 => x"65736829",
   643 => x"20617420",
   644 => x"30202867",
   645 => x"6f742030",
   646 => x"78256429",
   647 => x"0a000000",
   648 => x"42797465",
   649 => x"20636865",
   650 => x"636b2066",
   651 => x"61696c65",
   652 => x"64202862",
   653 => x"65666f72",
   654 => x"65206361",
   655 => x"63686520",
   656 => x"72656672",
   657 => x"65736829",
   658 => x"20617420",
   659 => x"33202867",
   660 => x"6f742030",
   661 => x"78256429",
   662 => x"0a000000",
   663 => x"42797465",
   664 => x"20636865",
   665 => x"636b2066",
   666 => x"61696c65",
   667 => x"64202861",
   668 => x"66746572",
   669 => x"20636163",
   670 => x"68652072",
   671 => x"65667265",
   672 => x"73682920",
   673 => x"61742030",
   674 => x"2028676f",
   675 => x"74203078",
   676 => x"2564290a",
   677 => x"00000000",
   678 => x"42797465",
   679 => x"20636865",
   680 => x"636b2066",
   681 => x"61696c65",
   682 => x"64202861",
   683 => x"66746572",
   684 => x"20636163",
   685 => x"68652072",
   686 => x"65667265",
   687 => x"73682920",
   688 => x"61742033",
   689 => x"2028676f",
   690 => x"74203078",
   691 => x"2564290a",
   692 => x"00000000",
   693 => x"43686563",
   694 => x"6b696e67",
   695 => x"206d656d",
   696 => x"6f727900",
   697 => x"30782564",
   698 => x"20676f6f",
   699 => x"64207265",
   700 => x"6164732c",
   701 => x"20000000",
   702 => x"4572726f",
   703 => x"72206174",
   704 => x"20307825",
   705 => x"642c2065",
   706 => x"78706563",
   707 => x"74656420",
   708 => x"30782564",
   709 => x"2c20676f",
   710 => x"74203078",
   711 => x"25640a00",
   712 => x"42616420",
   713 => x"64617461",
   714 => x"20666f75",
   715 => x"6e642061",
   716 => x"74203078",
   717 => x"25642028",
   718 => x"30782564",
   719 => x"290a0000",
   720 => x"53445241",
   721 => x"4d207369",
   722 => x"7a652028",
   723 => x"61737375",
   724 => x"6d696e67",
   725 => x"206e6f20",
   726 => x"61646472",
   727 => x"65737320",
   728 => x"6661756c",
   729 => x"74732920",
   730 => x"69732030",
   731 => x"78256420",
   732 => x"6d656761",
   733 => x"62797465",
   734 => x"730a0000",
   735 => x"416c6961",
   736 => x"73657320",
   737 => x"666f756e",
   738 => x"64206174",
   739 => x"20307825",
   740 => x"640a0000",
   741 => x"28416c69",
   742 => x"61736573",
   743 => x"2070726f",
   744 => x"6261626c",
   745 => x"79207369",
   746 => x"6d706c79",
   747 => x"20696e64",
   748 => x"69636174",
   749 => x"65207468",
   750 => x"61742052",
   751 => x"414d0a69",
   752 => x"7320736d",
   753 => x"616c6c65",
   754 => x"72207468",
   755 => x"616e2036",
   756 => x"34206d65",
   757 => x"67616279",
   758 => x"74657329",
   759 => x"0a000000",
   760 => x"46697273",
   761 => x"74207374",
   762 => x"61676520",
   763 => x"73616e69",
   764 => x"74792063",
   765 => x"6865636b",
   766 => x"20706173",
   767 => x"7365642e",
   768 => x"0a000000",
   769 => x"42797465",
   770 => x"20286471",
   771 => x"6d292063",
   772 => x"6865636b",
   773 => x"20706173",
   774 => x"7365640a",
   775 => x"00000000",
   776 => x"4c465352",
   777 => x"20636865",
   778 => x"636b2070",
   779 => x"61737365",
   780 => x"642e0a0a",
   781 => x"00000000",
   782 => x"41646472",
   783 => x"65737320",
   784 => x"63686563",
   785 => x"6b207061",
   786 => x"73736564",
   787 => x"2e0a0000",
	others => x"00000000"
);

begin

process (clk)
begin
	if (clk'event and clk = '1') then
		if (from_zpu.memAWriteEnable = '1') and (from_zpu.memBWriteEnable = '1') and (from_zpu.memAAddr=from_zpu.memBAddr) and (from_zpu.memAWrite/=from_zpu.memBWrite) then
			report "write collision" severity failure;
		end if;
	
		if (from_zpu.memAWriteEnable = '1') then
			ram(to_integer(unsigned(from_zpu.memAAddr(maxAddrBitBRAM downto 2)))) := from_zpu.memAWrite;
			to_zpu.memARead <= from_zpu.memAWrite;
		else
			to_zpu.memARead <= ram(to_integer(unsigned(from_zpu.memAAddr(maxAddrBitBRAM downto 2))));
		end if;
	end if;
end process;

process (clk)
begin
	if (clk'event and clk = '1') then
		if (from_zpu.memBWriteEnable = '1') then
			ram(to_integer(unsigned(from_zpu.memBAddr(maxAddrBitBRAM downto 2)))) := from_zpu.memBWrite;
			to_zpu.memBRead <= from_zpu.memBWrite;
		else
			to_zpu.memBRead <= ram(to_integer(unsigned(from_zpu.memBAddr(maxAddrBitBRAM downto 2))));
		end if;
	end if;
end process;


end arch;

