-- ZPU
--
-- Copyright 2004-2008 oharboe - �yvind Harboe - oyvind.harboe@zylin.com
-- Modified by Alastair M. Robinson for the ZPUFlex project.
--
-- The FreeBSD license
-- 
-- Redistribution and use in source and binary forms, with or without
-- modification, are permitted provided that the following conditions
-- are met:
-- 
-- 1. Redistributions of source code must retain the above copyright
--    notice, this list of conditions and the following disclaimer.
-- 2. Redistributions in binary form must reproduce the above
--    copyright notice, this list of conditions and the following
--    disclaimer in the documentation and/or other materials
--    provided with the distribution.
-- 
-- THIS SOFTWARE IS PROVIDED BY THE ZPU PROJECT ``AS IS'' AND ANY
-- EXPRESS OR IMPLIED WARRANTIES, INCLUDING, BUT NOT LIMITED TO,
-- THE IMPLIED WARRANTIES OF MERCHANTABILITY AND FITNESS FOR A
-- PARTICULAR PURPOSE ARE DISCLAIMED. IN NO EVENT SHALL THE
-- ZPU PROJECT OR CONTRIBUTORS BE LIABLE FOR ANY DIRECT,
-- INDIRECT, INCIDENTAL, SPECIAL, EXEMPLARY, OR CONSEQUENTIAL DAMAGES
-- (INCLUDING, BUT NOT LIMITED TO, PROCUREMENT OF SUBSTITUTE GOODS
-- OR SERVICES; LOSS OF USE, DATA, OR PROFITS; OR BUSINESS INTERRUPTION)
-- HOWEVER CAUSED AND ON ANY THEORY OF LIABILITY, WHETHER IN CONTRACT,
-- STRICT LIABILITY, OR TORT (INCLUDING NEGLIGENCE OR OTHERWISE)
-- ARISING IN ANY WAY OUT OF THE USE OF THIS SOFTWARE, EVEN IF
-- ADVISED OF THE POSSIBILITY OF SUCH DAMAGE.
-- 
-- The views and conclusions contained in the software and documentation
-- are those of the authors and should not be interpreted as representing
-- official policies, either expressed or implied, of the ZPU Project.

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;


library work;
use work.zpu_config.all;
use work.zpupkg.all;

entity SDBootstrap_ROM is
generic
	(
		maxAddrBit : integer := maxAddrBitBRAMLimit -- Specify your actual ROM size to save LEs and unnecessary block RAM usage.
	);
port (
	clk : in std_logic;
	areset : in std_logic := '0';
	from_zpu : in ZPU_ToROM;
	to_zpu : out ZPU_FromROM
);
end SDBootstrap_ROM;

architecture arch of SDBootstrap_ROM is

type ram_type is array(natural range 0 to ((2**(maxAddrBit+1))/4)-1) of std_logic_vector(wordSize-1 downto 0);

shared variable ram : ram_type :=
(
     0 => x"0ba08080",
     1 => x"ec040000",
     2 => x"00000000",
     3 => x"0ba08080",
     4 => x"880d8004",
     5 => x"a0808094",
     6 => x"0471fd06",
     7 => x"08728306",
     8 => x"09810582",
     9 => x"05832b2a",
    10 => x"83ffff06",
    11 => x"520471fc",
    12 => x"06087283",
    13 => x"06098105",
    14 => x"83051010",
    15 => x"102a81ff",
    16 => x"06520471",
    17 => x"fc06080b",
    18 => x"a0809ef0",
    19 => x"73830610",
    20 => x"10050806",
    21 => x"7381ff06",
    22 => x"73830609",
    23 => x"81058305",
    24 => x"1010102b",
    25 => x"0772fc06",
    26 => x"0c515104",
    27 => x"0284050b",
    28 => x"a0808088",
    29 => x"0ca08080",
    30 => x"940ba080",
    31 => x"8d9b0400",
    32 => x"0002c405",
    33 => x"0d0280c0",
    34 => x"0583ffe0",
    35 => x"e05b5680",
    36 => x"76708405",
    37 => x"5808715e",
    38 => x"5e577c70",
    39 => x"84055e08",
    40 => x"58805b77",
    41 => x"982a7888",
    42 => x"2b595372",
    43 => x"8838765e",
    44 => x"a08083aa",
    45 => x"047b802e",
    46 => x"81ca3880",
    47 => x"5c7280e4",
    48 => x"2e9f3872",
    49 => x"80e4268d",
    50 => x"387280e3",
    51 => x"2e80ee38",
    52 => x"a08082ca",
    53 => x"047280f3",
    54 => x"2e80cc38",
    55 => x"a08082ca",
    56 => x"04758417",
    57 => x"71087e5c",
    58 => x"56575287",
    59 => x"55739c2a",
    60 => x"74842b55",
    61 => x"5271802e",
    62 => x"83388159",
    63 => x"89722589",
    64 => x"38b71252",
    65 => x"a080828c",
    66 => x"04b01252",
    67 => x"78802e88",
    68 => x"387151a0",
    69 => x"8083b52d",
    70 => x"ff155574",
    71 => x"8025ce38",
    72 => x"8054a080",
    73 => x"82e00475",
    74 => x"84177108",
    75 => x"70545c57",
    76 => x"52a08083",
    77 => x"d92d7b54",
    78 => x"a08082e0",
    79 => x"04758417",
    80 => x"71085557",
    81 => x"52a08083",
    82 => x"9304a551",
    83 => x"a08083b5",
    84 => x"2d7251a0",
    85 => x"8083b52d",
    86 => x"821757a0",
    87 => x"80839d04",
    88 => x"73ff1555",
    89 => x"52807225",
    90 => x"b4387970",
    91 => x"81055ba0",
    92 => x"8080ae2d",
    93 => x"705253a0",
    94 => x"8083b52d",
    95 => x"811757a0",
    96 => x"8082e004",
    97 => x"72a52e09",
    98 => x"81068838",
    99 => x"815ca080",
   100 => x"839d0472",
   101 => x"51a08083",
   102 => x"b52d8117",
   103 => x"57811b5b",
   104 => x"837b25fd",
   105 => x"fe3872fd",
   106 => x"f1387d83",
   107 => x"ffe0800c",
   108 => x"02bc050d",
   109 => x"0402f805",
   110 => x"0d7352c0",
   111 => x"0870882a",
   112 => x"70810651",
   113 => x"51517080",
   114 => x"2ef13871",
   115 => x"c00c7183",
   116 => x"ffe0800c",
   117 => x"0288050d",
   118 => x"0402e805",
   119 => x"0d775574",
   120 => x"70840556",
   121 => x"08538054",
   122 => x"72982a73",
   123 => x"882b5452",
   124 => x"71802ea2",
   125 => x"38c00870",
   126 => x"882a7081",
   127 => x"06515151",
   128 => x"70802ef1",
   129 => x"3871c00c",
   130 => x"81168115",
   131 => x"55568374",
   132 => x"25d63871",
   133 => x"ca387583",
   134 => x"ffe0800c",
   135 => x"0298050d",
   136 => x"0402f405",
   137 => x"0d747671",
   138 => x"81ff06d4",
   139 => x"0c535383",
   140 => x"fff1a008",
   141 => x"85387189",
   142 => x"2b527198",
   143 => x"2ad40c71",
   144 => x"902a7081",
   145 => x"ff06d40c",
   146 => x"5171882a",
   147 => x"7081ff06",
   148 => x"d40c5171",
   149 => x"81ff06d4",
   150 => x"0c72902a",
   151 => x"7081ff06",
   152 => x"d40c51d4",
   153 => x"087081ff",
   154 => x"06515182",
   155 => x"b8bf5270",
   156 => x"81ff2e09",
   157 => x"81069438",
   158 => x"81ff0bd4",
   159 => x"0cd40870",
   160 => x"81ff06ff",
   161 => x"14545151",
   162 => x"71e53870",
   163 => x"83ffe080",
   164 => x"0c028c05",
   165 => x"0d0402fc",
   166 => x"050d81c7",
   167 => x"5181ff0b",
   168 => x"d40cff11",
   169 => x"51708025",
   170 => x"f4380284",
   171 => x"050d0402",
   172 => x"f0050da0",
   173 => x"8085962d",
   174 => x"819c9f53",
   175 => x"805287fc",
   176 => x"80f751a0",
   177 => x"8084a12d",
   178 => x"83ffe080",
   179 => x"085483ff",
   180 => x"e0800881",
   181 => x"2e098106",
   182 => x"ab3881ff",
   183 => x"0bd40c82",
   184 => x"0a52849c",
   185 => x"80e951a0",
   186 => x"8084a12d",
   187 => x"83ffe080",
   188 => x"088d3881",
   189 => x"ff0bd40c",
   190 => x"7353a080",
   191 => x"868b04a0",
   192 => x"8085962d",
   193 => x"ff135372",
   194 => x"ffb23872",
   195 => x"83ffe080",
   196 => x"0c029005",
   197 => x"0d0402f4",
   198 => x"050d81ff",
   199 => x"0bd40ca0",
   200 => x"809f8051",
   201 => x"a08083d9",
   202 => x"2d935380",
   203 => x"5287fc80",
   204 => x"c151a080",
   205 => x"84a12d83",
   206 => x"ffe08008",
   207 => x"8d3881ff",
   208 => x"0bd40c81",
   209 => x"53a08086",
   210 => x"d504a080",
   211 => x"85962dff",
   212 => x"135372d7",
   213 => x"387283ff",
   214 => x"e0800c02",
   215 => x"8c050d04",
   216 => x"02f0050d",
   217 => x"a0808596",
   218 => x"2d83aa52",
   219 => x"849c80c8",
   220 => x"51a08084",
   221 => x"a12d83ff",
   222 => x"e0800883",
   223 => x"ffe08008",
   224 => x"53a0809f",
   225 => x"8c5254a0",
   226 => x"8081812d",
   227 => x"73812e09",
   228 => x"81069038",
   229 => x"d8087083",
   230 => x"ffff0654",
   231 => x"547283aa",
   232 => x"2ea338a0",
   233 => x"8086962d",
   234 => x"a08087be",
   235 => x"048154a0",
   236 => x"8088f304",
   237 => x"a0809fa4",
   238 => x"51a08081",
   239 => x"812d8054",
   240 => x"a08088f3",
   241 => x"047352a0",
   242 => x"809fc051",
   243 => x"a0808181",
   244 => x"2d81ff0b",
   245 => x"d40cb153",
   246 => x"a08085af",
   247 => x"2d83ffe0",
   248 => x"8008802e",
   249 => x"80f43880",
   250 => x"5287fc80",
   251 => x"fa51a080",
   252 => x"84a12d83",
   253 => x"ffe08008",
   254 => x"80d03883",
   255 => x"ffe08008",
   256 => x"52a0809f",
   257 => x"d851a080",
   258 => x"81812d81",
   259 => x"ff0bd40c",
   260 => x"d40881ff",
   261 => x"067053a0",
   262 => x"809fe452",
   263 => x"54a08081",
   264 => x"812d81ff",
   265 => x"0bd40c81",
   266 => x"ff0bd40c",
   267 => x"81ff0bd4",
   268 => x"0c81ff0b",
   269 => x"d40c7386",
   270 => x"2a708106",
   271 => x"70565153",
   272 => x"72802eaf",
   273 => x"38a08087",
   274 => x"ad0483ff",
   275 => x"e0800852",
   276 => x"a0809fd8",
   277 => x"51a08081",
   278 => x"812d7282",
   279 => x"2efed538",
   280 => x"ff135372",
   281 => x"fef238a0",
   282 => x"809ff451",
   283 => x"a08083d9",
   284 => x"2d725473",
   285 => x"83ffe080",
   286 => x"0c029005",
   287 => x"0d0402f4",
   288 => x"050d810b",
   289 => x"83fff1a0",
   290 => x"0cd00870",
   291 => x"8f2a7081",
   292 => x"06515153",
   293 => x"72f33872",
   294 => x"d00ca080",
   295 => x"85962da0",
   296 => x"80a08c51",
   297 => x"a08083d9",
   298 => x"2dd00870",
   299 => x"8f2a7081",
   300 => x"06515153",
   301 => x"72f33881",
   302 => x"0bd00c87",
   303 => x"53805284",
   304 => x"d480c051",
   305 => x"a08084a1",
   306 => x"2d83ffe0",
   307 => x"8008812e",
   308 => x"09810687",
   309 => x"3883ffe0",
   310 => x"800853a0",
   311 => x"80a09c51",
   312 => x"a08083d9",
   313 => x"2d72822e",
   314 => x"09810692",
   315 => x"38a080a0",
   316 => x"b051a080",
   317 => x"83d92d80",
   318 => x"53a0808a",
   319 => x"ee04ff13",
   320 => x"5372ffb9",
   321 => x"38a080a0",
   322 => x"d051a080",
   323 => x"83d92da0",
   324 => x"8086e02d",
   325 => x"83ffe080",
   326 => x"0883fff1",
   327 => x"a00c83ff",
   328 => x"e0800880",
   329 => x"2e8b38a0",
   330 => x"80a0ec51",
   331 => x"a08083d9",
   332 => x"2da080a1",
   333 => x"8051a080",
   334 => x"83d92d81",
   335 => x"5287fc80",
   336 => x"d051a080",
   337 => x"84a12d81",
   338 => x"ff0bd40c",
   339 => x"d008708f",
   340 => x"2a708106",
   341 => x"51515372",
   342 => x"f33872d0",
   343 => x"0c81ff0b",
   344 => x"d40ca080",
   345 => x"a19051a0",
   346 => x"8083d92d",
   347 => x"81537283",
   348 => x"ffe0800c",
   349 => x"028c050d",
   350 => x"04800b83",
   351 => x"ffe0800c",
   352 => x"0402e005",
   353 => x"0d797b57",
   354 => x"57805881",
   355 => x"ff0bd40c",
   356 => x"d008708f",
   357 => x"2a708106",
   358 => x"51515473",
   359 => x"f3388281",
   360 => x"0bd00c81",
   361 => x"ff0bd40c",
   362 => x"765287fc",
   363 => x"80d151a0",
   364 => x"8084a12d",
   365 => x"80dbc6df",
   366 => x"5583ffe0",
   367 => x"8008802e",
   368 => x"983883ff",
   369 => x"e0800853",
   370 => x"7652a080",
   371 => x"a19c51a0",
   372 => x"8081812d",
   373 => x"a0808ca5",
   374 => x"0481ff0b",
   375 => x"d40cd408",
   376 => x"7081ff06",
   377 => x"51547381",
   378 => x"fe2e0981",
   379 => x"069b3880",
   380 => x"ff55d808",
   381 => x"76708405",
   382 => x"580cff15",
   383 => x"55748025",
   384 => x"f1388158",
   385 => x"a0808c8f",
   386 => x"04ff1555",
   387 => x"74cb3881",
   388 => x"ff0bd40c",
   389 => x"d008708f",
   390 => x"2a708106",
   391 => x"51515473",
   392 => x"f33873d0",
   393 => x"0c7783ff",
   394 => x"e0800c02",
   395 => x"a0050d04",
   396 => x"02f4050d",
   397 => x"7470882a",
   398 => x"83fe8006",
   399 => x"7072982a",
   400 => x"0772882b",
   401 => x"87fc8080",
   402 => x"0673982b",
   403 => x"81f00a06",
   404 => x"71730707",
   405 => x"83ffe080",
   406 => x"0c565153",
   407 => x"51028c05",
   408 => x"0d0402f8",
   409 => x"050d028e",
   410 => x"05a08080",
   411 => x"ae2d7498",
   412 => x"2b71902b",
   413 => x"0770902c",
   414 => x"83ffe080",
   415 => x"0c525202",
   416 => x"88050d04",
   417 => x"02f8050d",
   418 => x"7370902b",
   419 => x"71902a07",
   420 => x"83ffe080",
   421 => x"0c520288",
   422 => x"050d0402",
   423 => x"ec050d80",
   424 => x"0b870a0c",
   425 => x"a080a1bc",
   426 => x"51a08083",
   427 => x"d92da080",
   428 => x"88fe2d83",
   429 => x"ffe08008",
   430 => x"802e81ef",
   431 => x"38a080a1",
   432 => x"d451a080",
   433 => x"83d92da0",
   434 => x"8090892d",
   435 => x"83ffe1a0",
   436 => x"52a080a1",
   437 => x"ec51a080",
   438 => x"9c922d83",
   439 => x"ffe08008",
   440 => x"802e81c7",
   441 => x"3883ffe1",
   442 => x"a00ba080",
   443 => x"a1f85254",
   444 => x"a08083d9",
   445 => x"2d805573",
   446 => x"70810555",
   447 => x"a08080ae",
   448 => x"2d5372a0",
   449 => x"2e80de38",
   450 => x"72a32e81",
   451 => x"86387280",
   452 => x"c72e0981",
   453 => x"068b38a0",
   454 => x"80808c2d",
   455 => x"a0808ec1",
   456 => x"04728a2e",
   457 => x"0981068b",
   458 => x"38a08080",
   459 => x"942da080",
   460 => x"8ec10472",
   461 => x"80cc2e09",
   462 => x"81068638",
   463 => x"83ffe1a0",
   464 => x"547281df",
   465 => x"06f00570",
   466 => x"81ff0651",
   467 => x"53b87327",
   468 => x"8938ef13",
   469 => x"7081ff06",
   470 => x"51537484",
   471 => x"2b730755",
   472 => x"a0808df7",
   473 => x"0472a32e",
   474 => x"aa387370",
   475 => x"810555a0",
   476 => x"8080ae2d",
   477 => x"5372a02e",
   478 => x"f138ff14",
   479 => x"54800b8b",
   480 => x"15a08080",
   481 => x"c32d7452",
   482 => x"7351a080",
   483 => x"9c922d74",
   484 => x"870a0c73",
   485 => x"70810555",
   486 => x"a08080ae",
   487 => x"2d53728a",
   488 => x"2e098106",
   489 => x"ee38a080",
   490 => x"8df504a0",
   491 => x"80a28c51",
   492 => x"a08083d9",
   493 => x"2d800b83",
   494 => x"ffe0800c",
   495 => x"0294050d",
   496 => x"0402e805",
   497 => x"0d77797b",
   498 => x"58555580",
   499 => x"53727625",
   500 => x"ab387470",
   501 => x"810556a0",
   502 => x"8080ae2d",
   503 => x"74708105",
   504 => x"56a08080",
   505 => x"ae2d5252",
   506 => x"71712e88",
   507 => x"388151a0",
   508 => x"808ffe04",
   509 => x"811353a0",
   510 => x"808fcd04",
   511 => x"80517083",
   512 => x"ffe0800c",
   513 => x"0298050d",
   514 => x"0402d805",
   515 => x"0dff0b83",
   516 => x"fff5cc0c",
   517 => x"800b83ff",
   518 => x"f5e00ca0",
   519 => x"80a29851",
   520 => x"a08083d9",
   521 => x"2d83fff1",
   522 => x"b8528051",
   523 => x"a0808b81",
   524 => x"2d83ffe0",
   525 => x"80085483",
   526 => x"ffe08008",
   527 => x"9238a080",
   528 => x"a2a851a0",
   529 => x"8083d92d",
   530 => x"7355a080",
   531 => x"97ed04a0",
   532 => x"80a2bc51",
   533 => x"a08083d9",
   534 => x"2d805681",
   535 => x"0b83fff1",
   536 => x"ac0c8853",
   537 => x"a080a2d4",
   538 => x"5283fff1",
   539 => x"ee51a080",
   540 => x"8fc12d83",
   541 => x"ffe08008",
   542 => x"762e0981",
   543 => x"068b3883",
   544 => x"ffe08008",
   545 => x"83fff1ac",
   546 => x"0c8853a0",
   547 => x"80a2e052",
   548 => x"83fff28a",
   549 => x"51a0808f",
   550 => x"c12d83ff",
   551 => x"e080088b",
   552 => x"3883ffe0",
   553 => x"800883ff",
   554 => x"f1ac0c83",
   555 => x"fff1ac08",
   556 => x"52a080a2",
   557 => x"ec51a080",
   558 => x"81812d83",
   559 => x"fff1ac08",
   560 => x"802e81bb",
   561 => x"3883fff4",
   562 => x"fe0ba080",
   563 => x"80ae2d83",
   564 => x"fff4ff0b",
   565 => x"a08080ae",
   566 => x"2d71982b",
   567 => x"71902b07",
   568 => x"83fff580",
   569 => x"0ba08080",
   570 => x"ae2d7088",
   571 => x"2b720783",
   572 => x"fff5810b",
   573 => x"a08080ae",
   574 => x"2d710783",
   575 => x"fff5b60b",
   576 => x"a08080ae",
   577 => x"2d83fff5",
   578 => x"b70ba080",
   579 => x"80ae2d71",
   580 => x"882b0753",
   581 => x"5f54525a",
   582 => x"56575573",
   583 => x"81abaa2e",
   584 => x"09810693",
   585 => x"387551a0",
   586 => x"808cb02d",
   587 => x"83ffe080",
   588 => x"0856a080",
   589 => x"92cd0473",
   590 => x"82d4d52e",
   591 => x"9038a080",
   592 => x"a38051a0",
   593 => x"8083d92d",
   594 => x"a08094c5",
   595 => x"047552a0",
   596 => x"80a3a051",
   597 => x"a0808181",
   598 => x"2d83fff1",
   599 => x"b8527551",
   600 => x"a0808b81",
   601 => x"2d83ffe0",
   602 => x"80085583",
   603 => x"ffe08008",
   604 => x"802e84f9",
   605 => x"38a080a3",
   606 => x"b851a080",
   607 => x"83d92da0",
   608 => x"80a3e051",
   609 => x"a0808181",
   610 => x"2d8853a0",
   611 => x"80a2e052",
   612 => x"83fff28a",
   613 => x"51a0808f",
   614 => x"c12d83ff",
   615 => x"e080088d",
   616 => x"38810b83",
   617 => x"fff5e00c",
   618 => x"a08093d6",
   619 => x"048853a0",
   620 => x"80a2d452",
   621 => x"83fff1ee",
   622 => x"51a0808f",
   623 => x"c12d83ff",
   624 => x"e0800880",
   625 => x"2e9038a0",
   626 => x"80a3f851",
   627 => x"a0808181",
   628 => x"2da08094",
   629 => x"c50483ff",
   630 => x"f5b60ba0",
   631 => x"8080ae2d",
   632 => x"547380d5",
   633 => x"2e098106",
   634 => x"80db3883",
   635 => x"fff5b70b",
   636 => x"a08080ae",
   637 => x"2d547381",
   638 => x"aa2e0981",
   639 => x"0680c638",
   640 => x"800b83ff",
   641 => x"f1b80ba0",
   642 => x"8080ae2d",
   643 => x"56547481",
   644 => x"e92e8338",
   645 => x"81547481",
   646 => x"eb2e8c38",
   647 => x"80557375",
   648 => x"2e098106",
   649 => x"83c73883",
   650 => x"fff1c30b",
   651 => x"a08080ae",
   652 => x"2d557491",
   653 => x"3883fff1",
   654 => x"c40ba080",
   655 => x"80ae2d54",
   656 => x"73822e88",
   657 => x"388055a0",
   658 => x"8097ed04",
   659 => x"83fff1c5",
   660 => x"0ba08080",
   661 => x"ae2d7083",
   662 => x"fff5e80c",
   663 => x"ff0583ff",
   664 => x"f5dc0c83",
   665 => x"fff1c60b",
   666 => x"a08080ae",
   667 => x"2d83fff1",
   668 => x"c70ba080",
   669 => x"80ae2d58",
   670 => x"76057782",
   671 => x"80290570",
   672 => x"83fff5d0",
   673 => x"0c83fff1",
   674 => x"c80ba080",
   675 => x"80ae2d70",
   676 => x"83fff5c8",
   677 => x"0c83fff5",
   678 => x"e0085957",
   679 => x"5876802e",
   680 => x"81df3888",
   681 => x"53a080a2",
   682 => x"e05283ff",
   683 => x"f28a51a0",
   684 => x"808fc12d",
   685 => x"83ffe080",
   686 => x"0882b238",
   687 => x"83fff5e8",
   688 => x"0870842b",
   689 => x"83fff5b8",
   690 => x"0c7083ff",
   691 => x"f5e40c83",
   692 => x"fff1dd0b",
   693 => x"a08080ae",
   694 => x"2d83fff1",
   695 => x"dc0ba080",
   696 => x"80ae2d71",
   697 => x"82802905",
   698 => x"83fff1de",
   699 => x"0ba08080",
   700 => x"ae2d7084",
   701 => x"80802912",
   702 => x"83fff1df",
   703 => x"0ba08080",
   704 => x"ae2d7081",
   705 => x"800a2912",
   706 => x"7083fff1",
   707 => x"b00c83ff",
   708 => x"f5c80871",
   709 => x"2983fff5",
   710 => x"d0080570",
   711 => x"83fff5f0",
   712 => x"0c83fff1",
   713 => x"e50ba080",
   714 => x"80ae2d83",
   715 => x"fff1e40b",
   716 => x"a08080ae",
   717 => x"2d718280",
   718 => x"290583ff",
   719 => x"f1e60ba0",
   720 => x"8080ae2d",
   721 => x"70848080",
   722 => x"291283ff",
   723 => x"f1e70ba0",
   724 => x"8080ae2d",
   725 => x"70982b81",
   726 => x"f00a0672",
   727 => x"057083ff",
   728 => x"f1b40cfe",
   729 => x"117e2977",
   730 => x"0583fff5",
   731 => x"d80c5259",
   732 => x"5243545e",
   733 => x"51525952",
   734 => x"5d575957",
   735 => x"a08097eb",
   736 => x"0483fff1",
   737 => x"ca0ba080",
   738 => x"80ae2d83",
   739 => x"fff1c90b",
   740 => x"a08080ae",
   741 => x"2d718280",
   742 => x"29057083",
   743 => x"fff5b80c",
   744 => x"70a02983",
   745 => x"ff057089",
   746 => x"2a7083ff",
   747 => x"f5e40c83",
   748 => x"fff1cf0b",
   749 => x"a08080ae",
   750 => x"2d83fff1",
   751 => x"ce0ba080",
   752 => x"80ae2d71",
   753 => x"82802905",
   754 => x"7083fff1",
   755 => x"b00c7b71",
   756 => x"291e7083",
   757 => x"fff5d80c",
   758 => x"7d83fff1",
   759 => x"b40c7305",
   760 => x"83fff5f0",
   761 => x"0c555e51",
   762 => x"51555581",
   763 => x"557483ff",
   764 => x"e0800c02",
   765 => x"a8050d04",
   766 => x"02ec050d",
   767 => x"7670872c",
   768 => x"7180ff06",
   769 => x"57555383",
   770 => x"fff5e008",
   771 => x"8a387288",
   772 => x"2c7381ff",
   773 => x"06565473",
   774 => x"83fff5cc",
   775 => x"082ea838",
   776 => x"83fff1b8",
   777 => x"5283fff5",
   778 => x"d0081451",
   779 => x"a0808b81",
   780 => x"2d83ffe0",
   781 => x"80085383",
   782 => x"ffe08008",
   783 => x"802e80cb",
   784 => x"387383ff",
   785 => x"f5cc0c83",
   786 => x"fff5e008",
   787 => x"802ea038",
   788 => x"74842983",
   789 => x"fff1b805",
   790 => x"70085253",
   791 => x"a0808cb0",
   792 => x"2d83ffe0",
   793 => x"8008f00a",
   794 => x"0655a080",
   795 => x"99890474",
   796 => x"1083fff1",
   797 => x"b80570a0",
   798 => x"8080992d",
   799 => x"5253a080",
   800 => x"8ce22d83",
   801 => x"ffe08008",
   802 => x"55745372",
   803 => x"83ffe080",
   804 => x"0c029405",
   805 => x"0d0402cc",
   806 => x"050d7e60",
   807 => x"5e5b8056",
   808 => x"ff0b83ff",
   809 => x"f5cc0c83",
   810 => x"fff1b408",
   811 => x"83fff5d8",
   812 => x"08565783",
   813 => x"fff5e008",
   814 => x"762e8e38",
   815 => x"83fff5e8",
   816 => x"08842b59",
   817 => x"a08099d1",
   818 => x"0483fff5",
   819 => x"e408842b",
   820 => x"59805a79",
   821 => x"792781e1",
   822 => x"38798f06",
   823 => x"a0175754",
   824 => x"73a13874",
   825 => x"52a080a4",
   826 => x"9851a080",
   827 => x"81812d83",
   828 => x"fff1b852",
   829 => x"74518115",
   830 => x"55a0808b",
   831 => x"812d83ff",
   832 => x"f1b85680",
   833 => x"76a08080",
   834 => x"ae2d5558",
   835 => x"73782e83",
   836 => x"38815873",
   837 => x"81e52e81",
   838 => x"98388170",
   839 => x"7906555c",
   840 => x"73802e81",
   841 => x"8c388b16",
   842 => x"a08080ae",
   843 => x"2d980658",
   844 => x"7780fe38",
   845 => x"8b537c52",
   846 => x"7551a080",
   847 => x"8fc12d83",
   848 => x"ffe08008",
   849 => x"80eb389c",
   850 => x"160851a0",
   851 => x"808cb02d",
   852 => x"83ffe080",
   853 => x"08841c0c",
   854 => x"9a16a080",
   855 => x"80992d51",
   856 => x"a0808ce2",
   857 => x"2d83ffe0",
   858 => x"800883ff",
   859 => x"e0800855",
   860 => x"5583fff5",
   861 => x"e008802e",
   862 => x"9e389416",
   863 => x"a0808099",
   864 => x"2d51a080",
   865 => x"8ce22d83",
   866 => x"ffe08008",
   867 => x"902b83ff",
   868 => x"f00a0670",
   869 => x"16515473",
   870 => x"881c0c77",
   871 => x"7b0c7c52",
   872 => x"a080a4b8",
   873 => x"51a08081",
   874 => x"812d7b54",
   875 => x"a0809c87",
   876 => x"04811a5a",
   877 => x"a08099d3",
   878 => x"0483fff5",
   879 => x"e008802e",
   880 => x"80c33876",
   881 => x"51a08097",
   882 => x"f82d83ff",
   883 => x"e0800883",
   884 => x"ffe08008",
   885 => x"53a080a4",
   886 => x"cc5257a0",
   887 => x"8081812d",
   888 => x"7680ffff",
   889 => x"fff80654",
   890 => x"7380ffff",
   891 => x"fff82e95",
   892 => x"38fe1783",
   893 => x"fff5e808",
   894 => x"2983fff5",
   895 => x"f0080555",
   896 => x"a08099d1",
   897 => x"04805473",
   898 => x"83ffe080",
   899 => x"0c02b405",
   900 => x"0d0402e4",
   901 => x"050d787a",
   902 => x"715483ff",
   903 => x"f5bc5355",
   904 => x"55a08099",
   905 => x"962d83ff",
   906 => x"e0800881",
   907 => x"ff065372",
   908 => x"802e8183",
   909 => x"38a080a4",
   910 => x"e451a080",
   911 => x"83d92d83",
   912 => x"fff5c008",
   913 => x"83ff0589",
   914 => x"2a578070",
   915 => x"56567577",
   916 => x"25818038",
   917 => x"83fff5c4",
   918 => x"08fe0583",
   919 => x"fff5e808",
   920 => x"2983fff5",
   921 => x"f0081176",
   922 => x"83fff5dc",
   923 => x"08060575",
   924 => x"545253a0",
   925 => x"808b812d",
   926 => x"83ffe080",
   927 => x"08802e80",
   928 => x"c7388115",
   929 => x"7083fff5",
   930 => x"dc080654",
   931 => x"55729638",
   932 => x"83fff5c4",
   933 => x"0851a080",
   934 => x"97f82d83",
   935 => x"ffe08008",
   936 => x"83fff5c4",
   937 => x"0c848014",
   938 => x"81175754",
   939 => x"767624ff",
   940 => x"a338a080",
   941 => x"9dd30474",
   942 => x"52a080a5",
   943 => x"8051a080",
   944 => x"81812da0",
   945 => x"809dd504",
   946 => x"83ffe080",
   947 => x"0853a080",
   948 => x"9dd50481",
   949 => x"537283ff",
   950 => x"e0800c02",
   951 => x"9c050d04",
   952 => x"83ffe08c",
   953 => x"080283ff",
   954 => x"e08c0cff",
   955 => x"3d0d800b",
   956 => x"83ffe08c",
   957 => x"08fc050c",
   958 => x"83ffe08c",
   959 => x"08880508",
   960 => x"8106ff11",
   961 => x"70097083",
   962 => x"ffe08c08",
   963 => x"8c050806",
   964 => x"83ffe08c",
   965 => x"08fc0508",
   966 => x"1183ffe0",
   967 => x"8c08fc05",
   968 => x"0c83ffe0",
   969 => x"8c088805",
   970 => x"08812a83",
   971 => x"ffe08c08",
   972 => x"88050c83",
   973 => x"ffe08c08",
   974 => x"8c050810",
   975 => x"83ffe08c",
   976 => x"088c050c",
   977 => x"51515151",
   978 => x"83ffe08c",
   979 => x"08880508",
   980 => x"802e8438",
   981 => x"ffa23983",
   982 => x"ffe08c08",
   983 => x"fc050870",
   984 => x"83ffe080",
   985 => x"0c51833d",
   986 => x"0d83ffe0",
   987 => x"8c0c0400",
   988 => x"00ffffff",
   989 => x"ff00ffff",
   990 => x"ffff00ff",
   991 => x"ffffff00",
   992 => x"436d645f",
   993 => x"696e6974",
   994 => x"0a000000",
   995 => x"636d645f",
   996 => x"434d4438",
   997 => x"20726573",
   998 => x"706f6e73",
   999 => x"653a2025",
  1000 => x"640a0000",
  1001 => x"53444843",
  1002 => x"20496e69",
  1003 => x"7469616c",
  1004 => x"697a6174",
  1005 => x"696f6e20",
  1006 => x"6572726f",
  1007 => x"72210a00",
  1008 => x"434d4438",
  1009 => x"5f342072",
  1010 => x"6573706f",
  1011 => x"6e73653a",
  1012 => x"2025640a",
  1013 => x"00000000",
  1014 => x"434d4435",
  1015 => x"38202564",
  1016 => x"0a202000",
  1017 => x"434d4435",
  1018 => x"385f3220",
  1019 => x"25640a20",
  1020 => x"20000000",
  1021 => x"44657465",
  1022 => x"726d696e",
  1023 => x"65642053",
  1024 => x"44484320",
  1025 => x"73746174",
  1026 => x"75730a00",
  1027 => x"41637469",
  1028 => x"76617469",
  1029 => x"6e672043",
  1030 => x"530a0000",
  1031 => x"53656e74",
  1032 => x"20726573",
  1033 => x"65742063",
  1034 => x"6f6d6d61",
  1035 => x"6e640a00",
  1036 => x"53442063",
  1037 => x"61726420",
  1038 => x"696e6974",
  1039 => x"69616c69",
  1040 => x"7a617469",
  1041 => x"6f6e2065",
  1042 => x"72726f72",
  1043 => x"210a0000",
  1044 => x"43617264",
  1045 => x"20726573",
  1046 => x"706f6e64",
  1047 => x"65642074",
  1048 => x"6f207265",
  1049 => x"7365740a",
  1050 => x"00000000",
  1051 => x"53444843",
  1052 => x"20636172",
  1053 => x"64206465",
  1054 => x"74656374",
  1055 => x"65640a00",
  1056 => x"53656e64",
  1057 => x"696e6720",
  1058 => x"636d6431",
  1059 => x"360a0000",
  1060 => x"496e6974",
  1061 => x"20646f6e",
  1062 => x"650a0000",
  1063 => x"52656164",
  1064 => x"20636f6d",
  1065 => x"6d616e64",
  1066 => x"20666169",
  1067 => x"6c656420",
  1068 => x"61742025",
  1069 => x"64202825",
  1070 => x"64290a00",
  1071 => x"496e6974",
  1072 => x"69616c69",
  1073 => x"7a696e67",
  1074 => x"20534420",
  1075 => x"63617264",
  1076 => x"0a000000",
  1077 => x"48756e74",
  1078 => x"696e6720",
  1079 => x"666f7220",
  1080 => x"70617274",
  1081 => x"6974696f",
  1082 => x"6e0a0000",
  1083 => x"4d414e49",
  1084 => x"46455354",
  1085 => x"4d535400",
  1086 => x"50617273",
  1087 => x"696e6720",
  1088 => x"6d616e69",
  1089 => x"66657374",
  1090 => x"0a000000",
  1091 => x"52657475",
  1092 => x"726e696e",
  1093 => x"670a0000",
  1094 => x"52656164",
  1095 => x"696e6720",
  1096 => x"4d42520a",
  1097 => x"00000000",
  1098 => x"52656164",
  1099 => x"206f6620",
  1100 => x"4d425220",
  1101 => x"6661696c",
  1102 => x"65640a00",
  1103 => x"4d425220",
  1104 => x"73756363",
  1105 => x"65737366",
  1106 => x"756c6c79",
  1107 => x"20726561",
  1108 => x"640a0000",
  1109 => x"46415431",
  1110 => x"36202020",
  1111 => x"00000000",
  1112 => x"46415433",
  1113 => x"32202020",
  1114 => x"00000000",
  1115 => x"50617274",
  1116 => x"6974696f",
  1117 => x"6e636f75",
  1118 => x"6e742025",
  1119 => x"640a0000",
  1120 => x"4e6f2070",
  1121 => x"61727469",
  1122 => x"74696f6e",
  1123 => x"20736967",
  1124 => x"6e617475",
  1125 => x"72652066",
  1126 => x"6f756e64",
  1127 => x"0a000000",
  1128 => x"52656164",
  1129 => x"696e6720",
  1130 => x"626f6f74",
  1131 => x"20736563",
  1132 => x"746f7220",
  1133 => x"25640a00",
  1134 => x"52656164",
  1135 => x"20626f6f",
  1136 => x"74207365",
  1137 => x"63746f72",
  1138 => x"2066726f",
  1139 => x"6d206669",
  1140 => x"72737420",
  1141 => x"70617274",
  1142 => x"6974696f",
  1143 => x"6e0a0000",
  1144 => x"48756e74",
  1145 => x"696e6720",
  1146 => x"666f7220",
  1147 => x"66696c65",
  1148 => x"73797374",
  1149 => x"656d0a00",
  1150 => x"556e7375",
  1151 => x"70706f72",
  1152 => x"74656420",
  1153 => x"70617274",
  1154 => x"6974696f",
  1155 => x"6e207479",
  1156 => x"7065210d",
  1157 => x"00000000",
  1158 => x"52656164",
  1159 => x"696e6720",
  1160 => x"64697265",
  1161 => x"63746f72",
  1162 => x"79207365",
  1163 => x"63746f72",
  1164 => x"2025640a",
  1165 => x"00000000",
  1166 => x"66696c65",
  1167 => x"20222573",
  1168 => x"2220666f",
  1169 => x"756e640d",
  1170 => x"00000000",
  1171 => x"47657446",
  1172 => x"41544c69",
  1173 => x"6e6b2072",
  1174 => x"65747572",
  1175 => x"6e656420",
  1176 => x"25640a00",
  1177 => x"4f70656e",
  1178 => x"65642066",
  1179 => x"696c652c",
  1180 => x"206c6f61",
  1181 => x"64696e67",
  1182 => x"2e2e2e0a",
  1183 => x"00000000",
  1184 => x"43616e27",
  1185 => x"74206f70",
  1186 => x"656e2025",
  1187 => x"730a0000",
	others => x"00000000"
);

begin

process (clk)
begin
	if (clk'event and clk = '1') then
		if (from_zpu.memAWriteEnable = '1') and (from_zpu.memBWriteEnable = '1') and (from_zpu.memAAddr=from_zpu.memBAddr) and (from_zpu.memAWrite/=from_zpu.memBWrite) then
			report "write collision" severity failure;
		end if;
	
		if (from_zpu.memAWriteEnable = '1') then
			ram(to_integer(unsigned(from_zpu.memAAddr(maxAddrBit downto 2)))) := from_zpu.memAWrite;
			to_zpu.memARead <= from_zpu.memAWrite;
		else
			to_zpu.memARead <= ram(to_integer(unsigned(from_zpu.memAAddr(maxAddrBit downto 2))));
		end if;
	end if;
end process;

process (clk)
begin
	if (clk'event and clk = '1') then
		if (from_zpu.memBWriteEnable = '1') then
			ram(to_integer(unsigned(from_zpu.memBAddr(maxAddrBit downto 2)))) := from_zpu.memBWrite;
			to_zpu.memBRead <= from_zpu.memBWrite;
		else
			to_zpu.memBRead <= ram(to_integer(unsigned(from_zpu.memBAddr(maxAddrBit downto 2))));
		end if;
	end if;
end process;


end arch;

